
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_P4_adder_Nbit_blocks4 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_P4_adder_Nbit_blocks4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_95;

architecture SYN_ARCHBEH of nd2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_94;

architecture SYN_ARCHBEH of nd2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_93;

architecture SYN_ARCHBEH of nd2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_92;

architecture SYN_ARCHBEH of nd2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_91;

architecture SYN_ARCHBEH of nd2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_90;

architecture SYN_ARCHBEH of nd2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_89;

architecture SYN_ARCHBEH of nd2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_88;

architecture SYN_ARCHBEH of nd2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_87;

architecture SYN_ARCHBEH of nd2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_86;

architecture SYN_ARCHBEH of nd2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_85;

architecture SYN_ARCHBEH of nd2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_84;

architecture SYN_ARCHBEH of nd2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_83;

architecture SYN_ARCHBEH of nd2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_82;

architecture SYN_ARCHBEH of nd2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_81;

architecture SYN_ARCHBEH of nd2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_80;

architecture SYN_ARCHBEH of nd2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_79;

architecture SYN_ARCHBEH of nd2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_78;

architecture SYN_ARCHBEH of nd2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_77;

architecture SYN_ARCHBEH of nd2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_76;

architecture SYN_ARCHBEH of nd2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_75;

architecture SYN_ARCHBEH of nd2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_74;

architecture SYN_ARCHBEH of nd2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_73;

architecture SYN_ARCHBEH of nd2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_72;

architecture SYN_ARCHBEH of nd2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_71;

architecture SYN_ARCHBEH of nd2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_70;

architecture SYN_ARCHBEH of nd2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_69;

architecture SYN_ARCHBEH of nd2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_68;

architecture SYN_ARCHBEH of nd2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_67;

architecture SYN_ARCHBEH of nd2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_66;

architecture SYN_ARCHBEH of nd2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_65;

architecture SYN_ARCHBEH of nd2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_64;

architecture SYN_ARCHBEH of nd2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_63;

architecture SYN_ARCHBEH of nd2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_62;

architecture SYN_ARCHBEH of nd2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_61;

architecture SYN_ARCHBEH of nd2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_60;

architecture SYN_ARCHBEH of nd2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_59;

architecture SYN_ARCHBEH of nd2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_58;

architecture SYN_ARCHBEH of nd2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_57;

architecture SYN_ARCHBEH of nd2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_56;

architecture SYN_ARCHBEH of nd2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_55;

architecture SYN_ARCHBEH of nd2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_54;

architecture SYN_ARCHBEH of nd2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_53;

architecture SYN_ARCHBEH of nd2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_52;

architecture SYN_ARCHBEH of nd2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_51;

architecture SYN_ARCHBEH of nd2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_50;

architecture SYN_ARCHBEH of nd2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_49;

architecture SYN_ARCHBEH of nd2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_48;

architecture SYN_ARCHBEH of nd2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_47;

architecture SYN_ARCHBEH of nd2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_46;

architecture SYN_ARCHBEH of nd2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_45;

architecture SYN_ARCHBEH of nd2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_44;

architecture SYN_ARCHBEH of nd2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_43;

architecture SYN_ARCHBEH of nd2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_42;

architecture SYN_ARCHBEH of nd2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_41;

architecture SYN_ARCHBEH of nd2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_40;

architecture SYN_ARCHBEH of nd2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_39;

architecture SYN_ARCHBEH of nd2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_38;

architecture SYN_ARCHBEH of nd2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_37;

architecture SYN_ARCHBEH of nd2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_36;

architecture SYN_ARCHBEH of nd2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_35;

architecture SYN_ARCHBEH of nd2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_34;

architecture SYN_ARCHBEH of nd2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_33;

architecture SYN_ARCHBEH of nd2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_32;

architecture SYN_ARCHBEH of nd2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_31;

architecture SYN_ARCHBEH of nd2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_30;

architecture SYN_ARCHBEH of nd2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_29;

architecture SYN_ARCHBEH of nd2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_28;

architecture SYN_ARCHBEH of nd2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_27;

architecture SYN_ARCHBEH of nd2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_26;

architecture SYN_ARCHBEH of nd2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25;

architecture SYN_ARCHBEH of nd2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24;

architecture SYN_ARCHBEH of nd2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_23;

architecture SYN_ARCHBEH of nd2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_22;

architecture SYN_ARCHBEH of nd2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_21;

architecture SYN_ARCHBEH of nd2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_20;

architecture SYN_ARCHBEH of nd2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_19;

architecture SYN_ARCHBEH of nd2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_18;

architecture SYN_ARCHBEH of nd2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_17;

architecture SYN_ARCHBEH of nd2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_16;

architecture SYN_ARCHBEH of nd2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_15;

architecture SYN_ARCHBEH of nd2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_14;

architecture SYN_ARCHBEH of nd2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_13;

architecture SYN_ARCHBEH of nd2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_12;

architecture SYN_ARCHBEH of nd2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_11;

architecture SYN_ARCHBEH of nd2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_10;

architecture SYN_ARCHBEH of nd2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_9;

architecture SYN_ARCHBEH of nd2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_8;

architecture SYN_ARCHBEH of nd2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_7;

architecture SYN_ARCHBEH of nd2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_6;

architecture SYN_ARCHBEH of nd2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_5;

architecture SYN_ARCHBEH of nd2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_4;

architecture SYN_ARCHBEH of nd2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_3;

architecture SYN_ARCHBEH of nd2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_2;

architecture SYN_ARCHBEH of nd2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_1;

architecture SYN_ARCHBEH of nd2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_31 is

   port( A : in std_logic;  Y : out std_logic);

end iv_31;

architecture SYN_ARCHSTRUCT of iv_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_30 is

   port( A : in std_logic;  Y : out std_logic);

end iv_30;

architecture SYN_ARCHSTRUCT of iv_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_29 is

   port( A : in std_logic;  Y : out std_logic);

end iv_29;

architecture SYN_ARCHSTRUCT of iv_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_28 is

   port( A : in std_logic;  Y : out std_logic);

end iv_28;

architecture SYN_ARCHSTRUCT of iv_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_27 is

   port( A : in std_logic;  Y : out std_logic);

end iv_27;

architecture SYN_ARCHSTRUCT of iv_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_26 is

   port( A : in std_logic;  Y : out std_logic);

end iv_26;

architecture SYN_ARCHSTRUCT of iv_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_25 is

   port( A : in std_logic;  Y : out std_logic);

end iv_25;

architecture SYN_ARCHSTRUCT of iv_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_24 is

   port( A : in std_logic;  Y : out std_logic);

end iv_24;

architecture SYN_ARCHSTRUCT of iv_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_23 is

   port( A : in std_logic;  Y : out std_logic);

end iv_23;

architecture SYN_ARCHSTRUCT of iv_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_22 is

   port( A : in std_logic;  Y : out std_logic);

end iv_22;

architecture SYN_ARCHSTRUCT of iv_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_21 is

   port( A : in std_logic;  Y : out std_logic);

end iv_21;

architecture SYN_ARCHSTRUCT of iv_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_20 is

   port( A : in std_logic;  Y : out std_logic);

end iv_20;

architecture SYN_ARCHSTRUCT of iv_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_19 is

   port( A : in std_logic;  Y : out std_logic);

end iv_19;

architecture SYN_ARCHSTRUCT of iv_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_18 is

   port( A : in std_logic;  Y : out std_logic);

end iv_18;

architecture SYN_ARCHSTRUCT of iv_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_17 is

   port( A : in std_logic;  Y : out std_logic);

end iv_17;

architecture SYN_ARCHSTRUCT of iv_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_16 is

   port( A : in std_logic;  Y : out std_logic);

end iv_16;

architecture SYN_ARCHSTRUCT of iv_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_15 is

   port( A : in std_logic;  Y : out std_logic);

end iv_15;

architecture SYN_ARCHSTRUCT of iv_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_14 is

   port( A : in std_logic;  Y : out std_logic);

end iv_14;

architecture SYN_ARCHSTRUCT of iv_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_13 is

   port( A : in std_logic;  Y : out std_logic);

end iv_13;

architecture SYN_ARCHSTRUCT of iv_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_12 is

   port( A : in std_logic;  Y : out std_logic);

end iv_12;

architecture SYN_ARCHSTRUCT of iv_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_11 is

   port( A : in std_logic;  Y : out std_logic);

end iv_11;

architecture SYN_ARCHSTRUCT of iv_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_10 is

   port( A : in std_logic;  Y : out std_logic);

end iv_10;

architecture SYN_ARCHSTRUCT of iv_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_9 is

   port( A : in std_logic;  Y : out std_logic);

end iv_9;

architecture SYN_ARCHSTRUCT of iv_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_8 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8;

architecture SYN_ARCHSTRUCT of iv_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_7 is

   port( A : in std_logic;  Y : out std_logic);

end iv_7;

architecture SYN_ARCHSTRUCT of iv_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_6 is

   port( A : in std_logic;  Y : out std_logic);

end iv_6;

architecture SYN_ARCHSTRUCT of iv_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_5 is

   port( A : in std_logic;  Y : out std_logic);

end iv_5;

architecture SYN_ARCHSTRUCT of iv_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_4 is

   port( A : in std_logic;  Y : out std_logic);

end iv_4;

architecture SYN_ARCHSTRUCT of iv_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_3 is

   port( A : in std_logic;  Y : out std_logic);

end iv_3;

architecture SYN_ARCHSTRUCT of iv_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_2 is

   port( A : in std_logic;  Y : out std_logic);

end iv_2;

architecture SYN_ARCHSTRUCT of iv_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_1 is

   port( A : in std_logic;  Y : out std_logic);

end iv_1;

architecture SYN_ARCHSTRUCT of iv_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_31;

architecture SYN_ARCHSTRUCT of mux21_31 is

   component nd2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_31 port map( A => S, Y => n_S);
   NAND1 : nd2_93 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_92 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_91 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_30;

architecture SYN_ARCHSTRUCT of mux21_30 is

   component nd2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_30 port map( A => S, Y => n_S);
   NAND1 : nd2_90 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_89 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_88 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_29;

architecture SYN_ARCHSTRUCT of mux21_29 is

   component nd2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_29 port map( A => S, Y => n_S);
   NAND1 : nd2_87 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_86 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_85 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_28;

architecture SYN_ARCHSTRUCT of mux21_28 is

   component nd2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_28 port map( A => S, Y => n_S);
   NAND1 : nd2_84 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_83 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_82 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_27;

architecture SYN_ARCHSTRUCT of mux21_27 is

   component nd2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_27 port map( A => S, Y => n_S);
   NAND1 : nd2_81 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_80 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_79 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_26;

architecture SYN_ARCHSTRUCT of mux21_26 is

   component nd2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_26 port map( A => S, Y => n_S);
   NAND1 : nd2_78 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_77 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_76 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_25;

architecture SYN_ARCHSTRUCT of mux21_25 is

   component nd2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_25 port map( A => S, Y => n_S);
   NAND1 : nd2_75 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_74 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_73 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_24;

architecture SYN_ARCHSTRUCT of mux21_24 is

   component nd2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_24 port map( A => S, Y => n_S);
   NAND1 : nd2_72 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_71 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_70 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_23;

architecture SYN_ARCHSTRUCT of mux21_23 is

   component nd2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_23 port map( A => S, Y => n_S);
   NAND1 : nd2_69 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_68 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_67 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_22;

architecture SYN_ARCHSTRUCT of mux21_22 is

   component nd2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_22 port map( A => S, Y => n_S);
   NAND1 : nd2_66 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_65 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_64 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_21;

architecture SYN_ARCHSTRUCT of mux21_21 is

   component nd2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_21 port map( A => S, Y => n_S);
   NAND1 : nd2_63 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_62 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_61 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_20;

architecture SYN_ARCHSTRUCT of mux21_20 is

   component nd2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_20 port map( A => S, Y => n_S);
   NAND1 : nd2_60 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_59 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_58 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_19;

architecture SYN_ARCHSTRUCT of mux21_19 is

   component nd2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_19 port map( A => S, Y => n_S);
   NAND1 : nd2_57 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_56 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_55 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_18;

architecture SYN_ARCHSTRUCT of mux21_18 is

   component nd2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_18 port map( A => S, Y => n_S);
   NAND1 : nd2_54 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_53 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_52 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_17;

architecture SYN_ARCHSTRUCT of mux21_17 is

   component nd2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_17 port map( A => S, Y => n_S);
   NAND1 : nd2_51 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_50 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_49 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_16;

architecture SYN_ARCHSTRUCT of mux21_16 is

   component nd2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_16 port map( A => S, Y => n_S);
   NAND1 : nd2_48 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_47 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_46 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_15;

architecture SYN_ARCHSTRUCT of mux21_15 is

   component nd2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_15 port map( A => S, Y => n_S);
   NAND1 : nd2_45 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_44 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_43 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_14;

architecture SYN_ARCHSTRUCT of mux21_14 is

   component nd2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_14 port map( A => S, Y => n_S);
   NAND1 : nd2_42 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_41 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_40 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_13;

architecture SYN_ARCHSTRUCT of mux21_13 is

   component nd2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_13 port map( A => S, Y => n_S);
   NAND1 : nd2_39 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_38 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_37 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_12;

architecture SYN_ARCHSTRUCT of mux21_12 is

   component nd2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_12 port map( A => S, Y => n_S);
   NAND1 : nd2_36 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_35 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_34 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_11;

architecture SYN_ARCHSTRUCT of mux21_11 is

   component nd2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_11 port map( A => S, Y => n_S);
   NAND1 : nd2_33 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_32 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_31 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_10;

architecture SYN_ARCHSTRUCT of mux21_10 is

   component nd2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_10 port map( A => S, Y => n_S);
   NAND1 : nd2_30 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_29 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_28 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_9;

architecture SYN_ARCHSTRUCT of mux21_9 is

   component nd2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_9 port map( A => S, Y => n_S);
   NAND1 : nd2_27 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_26 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8;

architecture SYN_ARCHSTRUCT of mux21_8 is

   component nd2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8 port map( A => S, Y => n_S);
   NAND1 : nd2_24 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_23 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_22 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_7;

architecture SYN_ARCHSTRUCT of mux21_7 is

   component nd2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_7 port map( A => S, Y => n_S);
   NAND1 : nd2_21 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_20 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_19 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_6;

architecture SYN_ARCHSTRUCT of mux21_6 is

   component nd2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_6 port map( A => S, Y => n_S);
   NAND1 : nd2_18 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_17 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_16 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_5;

architecture SYN_ARCHSTRUCT of mux21_5 is

   component nd2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_5 port map( A => S, Y => n_S);
   NAND1 : nd2_15 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_14 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_13 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_4;

architecture SYN_ARCHSTRUCT of mux21_4 is

   component nd2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_4 port map( A => S, Y => n_S);
   NAND1 : nd2_12 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_11 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_10 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_3;

architecture SYN_ARCHSTRUCT of mux21_3 is

   component nd2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_3 port map( A => S, Y => n_S);
   NAND1 : nd2_9 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_8 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_7 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_2;

architecture SYN_ARCHSTRUCT of mux21_2 is

   component nd2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_2 port map( A => S, Y => n_S);
   NAND1 : nd2_6 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_5 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_4 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_1;

architecture SYN_ARCHSTRUCT of mux21_1 is

   component nd2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_1 port map( A => S, Y => n_S);
   NAND1 : nd2_3 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_2 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_1 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_ARCHBEH of FA_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_ARCHBEH of FA_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_ARCHBEH of FA_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_ARCHBEH of FA_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_ARCHBEH of FA_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_ARCHBEH of FA_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_ARCHBEH of FA_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_ARCHBEH of FA_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_ARCHBEH of FA_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_ARCHBEH of FA_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_ARCHBEH of FA_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_ARCHBEH of FA_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_ARCHBEH of FA_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_ARCHBEH of FA_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_ARCHBEH of FA_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_ARCHBEH of FA_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_ARCHBEH of FA_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_ARCHBEH of FA_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_ARCHBEH of FA_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_ARCHBEH of FA_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_ARCHBEH of FA_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_ARCHBEH of FA_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_ARCHBEH of FA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_ARCHBEH of FA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_ARCHBEH of FA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_ARCHBEH of FA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_ARCHBEH of FA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_ARCHBEH of FA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_ARCHBEH of FA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_ARCHBEH of FA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_ARCHBEH of FA_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_ARCHBEH of FA_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_ARCHBEH of FA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_ARCHBEH of FA_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_ARCHBEH of FA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_ARCHBEH of FA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_ARCHBEH of FA_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_ARCHBEH of FA_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_ARCHBEH of FA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_ARCHBEH of FA_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_ARCHBEH of FA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_ARCHBEH of FA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_ARCHBEH of FA_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_ARCHBEH of FA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_ARCHBEH of FA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_ARCHBEH of FA_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_ARCHBEH of FA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_ARCHBEH of FA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_ARCHBEH of FA_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_ARCHBEH of FA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_ARCHBEH of FA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_ARCHBEH of FA_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_ARCHBEH of FA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_ARCHBEH of FA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_ARCHBEH of FA_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_ARCHBEH of FA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_ARCHBEH of FA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_ARCHBEH of FA_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_ARCHBEH of FA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_ARCHBEH of FA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_ARCHBEH of FA_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_ARCHBEH of FA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_ARCHBEH of FA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity muxN1_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_7;

architecture SYN_ARCHSTRUCT of muxN1_N4_7 is

   component mux21_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_28 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_27 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_26 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_25 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity muxN1_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_6;

architecture SYN_ARCHSTRUCT of muxN1_N4_6 is

   component mux21_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_24 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_23 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_22 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_21 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity muxN1_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_5;

architecture SYN_ARCHSTRUCT of muxN1_N4_5 is

   component mux21_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_20 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_19 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_18 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_17 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity muxN1_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_4;

architecture SYN_ARCHSTRUCT of muxN1_N4_4 is

   component mux21_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_16 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_15 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_14 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_13 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity muxN1_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_3;

architecture SYN_ARCHSTRUCT of muxN1_N4_3 is

   component mux21_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_12 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_11 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_10 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_9 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity muxN1_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_2;

architecture SYN_ARCHSTRUCT of muxN1_N4_2 is

   component mux21_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_7 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_6 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_5 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity muxN1_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_1;

architecture SYN_ARCHSTRUCT of muxN1_N4_1 is

   component mux21_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_4 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_3 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_2 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_1 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_15;

architecture SYN_ARCHSTRUCT of RCA_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_14;

architecture SYN_ARCHSTRUCT of RCA_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_13;

architecture SYN_ARCHSTRUCT of RCA_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_12;

architecture SYN_ARCHSTRUCT of RCA_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_11;

architecture SYN_ARCHSTRUCT of RCA_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_10;

architecture SYN_ARCHSTRUCT of RCA_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_9;

architecture SYN_ARCHSTRUCT of RCA_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_8;

architecture SYN_ARCHSTRUCT of RCA_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_7;

architecture SYN_ARCHSTRUCT of RCA_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_6;

architecture SYN_ARCHSTRUCT of RCA_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_5;

architecture SYN_ARCHSTRUCT of RCA_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_4;

architecture SYN_ARCHSTRUCT of RCA_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_3;

architecture SYN_ARCHSTRUCT of RCA_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_2;

architecture SYN_ARCHSTRUCT of RCA_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_1;

architecture SYN_ARCHSTRUCT of RCA_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_26 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_26;

architecture SYN_ARCHDATAFLOW of pg_block_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_25 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_25;

architecture SYN_ARCHDATAFLOW of pg_block_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_24 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_24;

architecture SYN_ARCHDATAFLOW of pg_block_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_23 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_23;

architecture SYN_ARCHDATAFLOW of pg_block_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_22 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_22;

architecture SYN_ARCHDATAFLOW of pg_block_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_21 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_21;

architecture SYN_ARCHDATAFLOW of pg_block_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_20 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_20;

architecture SYN_ARCHDATAFLOW of pg_block_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_19 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_19;

architecture SYN_ARCHDATAFLOW of pg_block_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_18 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_18;

architecture SYN_ARCHDATAFLOW of pg_block_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_17 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_17;

architecture SYN_ARCHDATAFLOW of pg_block_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_16 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_16;

architecture SYN_ARCHDATAFLOW of pg_block_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_15 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_15;

architecture SYN_ARCHDATAFLOW of pg_block_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_14 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_14;

architecture SYN_ARCHDATAFLOW of pg_block_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_13 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_13;

architecture SYN_ARCHDATAFLOW of pg_block_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_12 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_12;

architecture SYN_ARCHDATAFLOW of pg_block_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_11 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_11;

architecture SYN_ARCHDATAFLOW of pg_block_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_10 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_10;

architecture SYN_ARCHDATAFLOW of pg_block_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_9 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_9;

architecture SYN_ARCHDATAFLOW of pg_block_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_8 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_8;

architecture SYN_ARCHDATAFLOW of pg_block_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_7 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_7;

architecture SYN_ARCHDATAFLOW of pg_block_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_6 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_6;

architecture SYN_ARCHDATAFLOW of pg_block_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_5 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_5;

architecture SYN_ARCHDATAFLOW of pg_block_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_4 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_4;

architecture SYN_ARCHDATAFLOW of pg_block_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_3 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_3;

architecture SYN_ARCHDATAFLOW of pg_block_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_2 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_2;

architecture SYN_ARCHDATAFLOW of pg_block_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_1 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_1;

architecture SYN_ARCHDATAFLOW of pg_block_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity g_block_8 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_8;

architecture SYN_ARCHDATAFLOW of g_block_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity g_block_7 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_7;

architecture SYN_ARCHDATAFLOW of g_block_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity g_block_6 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_6;

architecture SYN_ARCHDATAFLOW of g_block_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity g_block_5 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_5;

architecture SYN_ARCHDATAFLOW of g_block_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity g_block_4 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_4;

architecture SYN_ARCHDATAFLOW of g_block_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity g_block_3 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_3;

architecture SYN_ARCHDATAFLOW of g_block_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity g_block_2 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_2;

architecture SYN_ARCHDATAFLOW of g_block_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity g_block_1 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_1;

architecture SYN_ARCHDATAFLOW of g_block_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_select_block_N4_7 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_7;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_7 is

   component muxN1_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1000, n_1001 : 
      std_logic;

begin
   
   RCA1 : RCA_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1000);
   RCA2 : RCA_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S2_3_port, 
                           S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1001);
   MUX : muxN1_N4_7 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_select_block_N4_6 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_6;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_6 is

   component muxN1_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1002, n_1003 : 
      std_logic;

begin
   
   RCA1 : RCA_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1002);
   RCA2 : RCA_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S2_3_port, 
                           S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1003);
   MUX : muxN1_N4_6 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_select_block_N4_5 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_5;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_5 is

   component muxN1_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1004, n_1005 : 
      std_logic;

begin
   
   RCA1 : RCA_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1004);
   RCA2 : RCA_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S2_3_port, 
                           S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1005);
   MUX : muxN1_N4_5 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_select_block_N4_4 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_4;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_4 is

   component muxN1_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1006, n_1007 : 
      std_logic;

begin
   
   RCA1 : RCA_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1006);
   RCA2 : RCA_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S2_3_port, 
                           S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1007);
   MUX : muxN1_N4_4 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_select_block_N4_3 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_3;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_3 is

   component muxN1_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1008, n_1009 : 
      std_logic;

begin
   
   RCA1 : RCA_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1008);
   RCA2 : RCA_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S2_3_port, 
                           S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1009);
   MUX : muxN1_N4_3 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_select_block_N4_2 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_2;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_2 is

   component muxN1_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1010, n_1011 : 
      std_logic;

begin
   
   RCA1 : RCA_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1010);
   RCA2 : RCA_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S2_3_port, 
                           S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1011);
   MUX : muxN1_N4_2 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_select_block_N4_1 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_1;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_1 is

   component muxN1_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1012, n_1013 : 
      std_logic;

begin
   
   RCA1 : RCA_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1012);
   RCA2 : RCA_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S2_3_port, 
                           S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1013);
   MUX : muxN1_N4_1 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity nd2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_0;

architecture SYN_ARCHBEH of nd2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity iv_0 is

   port( A : in std_logic;  Y : out std_logic);

end iv_0;

architecture SYN_ARCHSTRUCT of iv_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity mux21_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_0;

architecture SYN_ARCHSTRUCT of mux21_0 is

   component nd2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_0 port map( A => S, Y => n_S);
   NAND1 : nd2_0 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_95 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_94 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_ARCHBEH of FA_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity muxN1_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_0;

architecture SYN_ARCHSTRUCT of muxN1_N4_0 is

   component mux21_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_0 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_31 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_30 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_29 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity RCA_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_0;

architecture SYN_ARCHSTRUCT of RCA_N4_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_block_0 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_0;

architecture SYN_ARCHDATAFLOW of pg_block_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);
   U2 : INV_X1 port map( A => n1, ZN => G_i_j);
   U3 : AOI21_X1 port map( B1 => G_kmin1_j, B2 => P_i_k, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity g_block_0 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_0;

architecture SYN_ARCHDATAFLOW of g_block_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_select_block_N4_0 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_0;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_0 is

   component muxN1_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1014, n_1015 : 
      std_logic;

begin
   
   RCA1 : RCA_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => S1_3_port, 
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1014);
   RCA2 : RCA_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) =>
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => S2_3_port, 
                           S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1015);
   MUX : muxN1_N4_0 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_generator_sparse_tree_N32_carry_range4 is

   port( P, G : in std_logic_vector (31 downto 0);  Cin : in std_logic;  C : 
         out std_logic_vector (8 downto 0));

end carry_generator_sparse_tree_N32_carry_range4;

architecture SYN_ARCHSTRUCT of carry_generator_sparse_tree_N32_carry_range4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component g_block_1
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component g_block_2
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component g_block_3
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component g_block_4
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_1
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_2
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_5
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component g_block_6
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_3
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_4
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_5
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_7
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_6
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_7
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_8
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_9
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_10
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_11
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_12
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_8
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_13
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_14
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_15
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_16
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_17
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_18
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_19
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_20
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_21
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_22
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_23
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_24
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_25
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_26
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_0
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_0
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   signal C_8_port, C_7_port, C_6_port, C_5_port, C_4_port, C_3_port, C_2_port,
      C_1_port, Gmat_16_15_port, Gmat_16_13_port, Gmat_16_9_port, 
      Gmat_14_13_port, Gmat_12_11_port, Gmat_12_9_port, Gmat_10_9_port, 
      Gmat_8_7_port, Gmat_8_5_port, Gmat_6_5_port, Gmat_4_3_port, Gmat_2_1_port
      , Pmat_16_15_port, Pmat_16_13_port, Pmat_16_9_port, Pmat_14_13_port, 
      Pmat_12_11_port, Pmat_12_9_port, Pmat_10_9_port, Pmat_8_7_port, 
      Pmat_8_5_port, Pmat_6_5_port, Pmat_4_3_port, Pmat_32_31_port, 
      Pmat_32_29_port, Pmat_32_25_port, Pmat_32_17_port, Pmat_30_29_port, 
      Pmat_28_27_port, Pmat_28_25_port, Pmat_28_17_port, Pmat_26_25_port, 
      Pmat_24_23_port, Pmat_24_21_port, Pmat_24_17_port, Pmat_22_21_port, 
      Pmat_20_19_port, Pmat_20_17_port, Pmat_18_17_port, Gmat_32_31_port, 
      Gmat_32_29_port, Gmat_32_25_port, Gmat_32_17_port, Gmat_30_29_port, 
      Gmat_28_27_port, Gmat_28_25_port, Gmat_28_17_port, Gmat_26_25_port, 
      Gmat_24_23_port, Gmat_24_21_port, Gmat_24_17_port, Gmat_22_21_port, 
      Gmat_20_19_port, Gmat_20_17_port, Gmat_18_17_port, n1, n2 : std_logic;

begin
   C <= ( C_8_port, C_7_port, C_6_port, C_5_port, C_4_port, C_3_port, C_2_port,
      C_1_port, Cin );
   
   first_G_1_2 : g_block_0 port map( G_i_k => G(1), G_kmin1_j => n1, P_i_k => 
                           P(1), G_i_j => Gmat_2_1_port);
   FRST_PG_1_4 : pg_block_0 port map( G_i_k => G(3), G_kmin1_j => G(2), P_i_k 
                           => P(3), P_kmin1_j => P(2), P_i_j => Pmat_4_3_port, 
                           G_i_j => Gmat_4_3_port);
   FRST_PG_1_6 : pg_block_26 port map( G_i_k => G(5), G_kmin1_j => G(4), P_i_k 
                           => P(5), P_kmin1_j => P(4), P_i_j => Pmat_6_5_port, 
                           G_i_j => Gmat_6_5_port);
   FRST_PG_1_8 : pg_block_25 port map( G_i_k => G(7), G_kmin1_j => G(6), P_i_k 
                           => P(7), P_kmin1_j => P(6), P_i_j => Pmat_8_7_port, 
                           G_i_j => Gmat_8_7_port);
   FRST_PG_1_10 : pg_block_24 port map( G_i_k => G(9), G_kmin1_j => G(8), P_i_k
                           => P(9), P_kmin1_j => P(8), P_i_j => Pmat_10_9_port,
                           G_i_j => Gmat_10_9_port);
   FRST_PG_1_12 : pg_block_23 port map( G_i_k => G(11), G_kmin1_j => G(10), 
                           P_i_k => P(11), P_kmin1_j => P(10), P_i_j => 
                           Pmat_12_11_port, G_i_j => Gmat_12_11_port);
   FRST_PG_1_14 : pg_block_22 port map( G_i_k => G(13), G_kmin1_j => G(12), 
                           P_i_k => P(13), P_kmin1_j => P(12), P_i_j => 
                           Pmat_14_13_port, G_i_j => Gmat_14_13_port);
   FRST_PG_1_16 : pg_block_21 port map( G_i_k => G(15), G_kmin1_j => G(14), 
                           P_i_k => P(15), P_kmin1_j => P(14), P_i_j => 
                           Pmat_16_15_port, G_i_j => Gmat_16_15_port);
   FRST_PG_1_18 : pg_block_20 port map( G_i_k => G(17), G_kmin1_j => G(16), 
                           P_i_k => P(17), P_kmin1_j => P(16), P_i_j => 
                           Pmat_18_17_port, G_i_j => Gmat_18_17_port);
   FRST_PG_1_20 : pg_block_19 port map( G_i_k => G(19), G_kmin1_j => G(18), 
                           P_i_k => P(19), P_kmin1_j => P(18), P_i_j => 
                           Pmat_20_19_port, G_i_j => Gmat_20_19_port);
   FRST_PG_1_22 : pg_block_18 port map( G_i_k => G(21), G_kmin1_j => G(20), 
                           P_i_k => P(21), P_kmin1_j => P(20), P_i_j => 
                           Pmat_22_21_port, G_i_j => Gmat_22_21_port);
   FRST_PG_1_24 : pg_block_17 port map( G_i_k => G(23), G_kmin1_j => G(22), 
                           P_i_k => P(23), P_kmin1_j => P(22), P_i_j => 
                           Pmat_24_23_port, G_i_j => Gmat_24_23_port);
   FRST_PG_1_26 : pg_block_16 port map( G_i_k => G(25), G_kmin1_j => G(24), 
                           P_i_k => P(25), P_kmin1_j => P(24), P_i_j => 
                           Pmat_26_25_port, G_i_j => Gmat_26_25_port);
   FRST_PG_1_28 : pg_block_15 port map( G_i_k => G(27), G_kmin1_j => G(26), 
                           P_i_k => P(27), P_kmin1_j => P(26), P_i_j => 
                           Pmat_28_27_port, G_i_j => Gmat_28_27_port);
   FRST_PG_1_30 : pg_block_14 port map( G_i_k => G(29), G_kmin1_j => G(28), 
                           P_i_k => P(29), P_kmin1_j => P(28), P_i_j => 
                           Pmat_30_29_port, G_i_j => Gmat_30_29_port);
   FRST_PG_1_32 : pg_block_13 port map( G_i_k => G(31), G_kmin1_j => G(30), 
                           P_i_k => P(31), P_kmin1_j => P(30), P_i_j => 
                           Pmat_32_31_port, G_i_j => Gmat_32_31_port);
   first_G_2_4 : g_block_8 port map( G_i_k => Gmat_4_3_port, G_kmin1_j => 
                           Gmat_2_1_port, P_i_k => Pmat_4_3_port, G_i_j => 
                           C_1_port);
   FRST_PG_2_8 : pg_block_12 port map( G_i_k => Gmat_8_7_port, G_kmin1_j => 
                           Gmat_6_5_port, P_i_k => Pmat_8_7_port, P_kmin1_j => 
                           Pmat_6_5_port, P_i_j => Pmat_8_5_port, G_i_j => 
                           Gmat_8_5_port);
   FRST_PG_2_12 : pg_block_11 port map( G_i_k => Gmat_12_11_port, G_kmin1_j => 
                           Gmat_10_9_port, P_i_k => Pmat_12_11_port, P_kmin1_j 
                           => Pmat_10_9_port, P_i_j => Pmat_12_9_port, G_i_j =>
                           Gmat_12_9_port);
   FRST_PG_2_16 : pg_block_10 port map( G_i_k => Gmat_16_15_port, G_kmin1_j => 
                           Gmat_14_13_port, P_i_k => Pmat_16_15_port, P_kmin1_j
                           => Pmat_14_13_port, P_i_j => Pmat_16_13_port, G_i_j 
                           => Gmat_16_13_port);
   FRST_PG_2_20 : pg_block_9 port map( G_i_k => Gmat_20_19_port, G_kmin1_j => 
                           Gmat_18_17_port, P_i_k => Pmat_20_19_port, P_kmin1_j
                           => Pmat_18_17_port, P_i_j => Pmat_20_17_port, G_i_j 
                           => Gmat_20_17_port);
   FRST_PG_2_24 : pg_block_8 port map( G_i_k => Gmat_24_23_port, G_kmin1_j => 
                           Gmat_22_21_port, P_i_k => Pmat_24_23_port, P_kmin1_j
                           => Pmat_22_21_port, P_i_j => Pmat_24_21_port, G_i_j 
                           => Gmat_24_21_port);
   FRST_PG_2_28 : pg_block_7 port map( G_i_k => Gmat_28_27_port, G_kmin1_j => 
                           Gmat_26_25_port, P_i_k => Pmat_28_27_port, P_kmin1_j
                           => Pmat_26_25_port, P_i_j => Pmat_28_25_port, G_i_j 
                           => Gmat_28_25_port);
   FRST_PG_2_32 : pg_block_6 port map( G_i_k => Gmat_32_31_port, G_kmin1_j => 
                           Gmat_30_29_port, P_i_k => Pmat_32_31_port, P_kmin1_j
                           => Pmat_30_29_port, P_i_j => Pmat_32_29_port, G_i_j 
                           => Gmat_32_29_port);
   G_L2_0_4_8 : g_block_7 port map( G_i_k => Gmat_8_5_port, G_kmin1_j => 
                           C_1_port, P_i_k => Pmat_8_5_port, G_i_j => C_2_port)
                           ;
   PG_L2_0_12_16 : pg_block_5 port map( G_i_k => Gmat_16_13_port, G_kmin1_j => 
                           Gmat_12_9_port, P_i_k => Pmat_16_13_port, P_kmin1_j 
                           => Pmat_12_9_port, P_i_j => Pmat_16_9_port, G_i_j =>
                           Gmat_16_9_port);
   PG_L2_0_20_24 : pg_block_4 port map( G_i_k => Gmat_24_21_port, G_kmin1_j => 
                           Gmat_20_17_port, P_i_k => Pmat_24_21_port, P_kmin1_j
                           => Pmat_20_17_port, P_i_j => Pmat_24_17_port, G_i_j 
                           => Gmat_24_17_port);
   PG_L2_0_28_32 : pg_block_3 port map( G_i_k => Gmat_32_29_port, G_kmin1_j => 
                           Gmat_28_25_port, P_i_k => Pmat_32_29_port, P_kmin1_j
                           => Pmat_28_25_port, P_i_j => Pmat_32_25_port, G_i_j 
                           => Gmat_32_25_port);
   G_L2_1_8_12 : g_block_6 port map( G_i_k => Gmat_12_9_port, G_kmin1_j => 
                           C_2_port, P_i_k => Pmat_12_9_port, G_i_j => C_3_port
                           );
   G_L2_1_8_16 : g_block_5 port map( G_i_k => Gmat_16_9_port, G_kmin1_j => 
                           C_2_port, P_i_k => Pmat_16_9_port, G_i_j => C_4_port
                           );
   PG_L2_1_24_28 : pg_block_2 port map( G_i_k => Gmat_28_25_port, G_kmin1_j => 
                           Gmat_24_17_port, P_i_k => Pmat_28_25_port, P_kmin1_j
                           => Pmat_24_17_port, P_i_j => Pmat_28_17_port, G_i_j 
                           => Gmat_28_17_port);
   PG_L2_1_24_32 : pg_block_1 port map( G_i_k => Gmat_32_25_port, G_kmin1_j => 
                           Gmat_24_17_port, P_i_k => Pmat_32_25_port, P_kmin1_j
                           => Pmat_24_17_port, P_i_j => Pmat_32_17_port, G_i_j 
                           => Gmat_32_17_port);
   G_L2_2_16_20 : g_block_4 port map( G_i_k => Gmat_20_17_port, G_kmin1_j => 
                           C_4_port, P_i_k => Pmat_20_17_port, G_i_j => 
                           C_5_port);
   G_L2_2_16_24 : g_block_3 port map( G_i_k => Gmat_24_17_port, G_kmin1_j => 
                           C_4_port, P_i_k => Pmat_24_17_port, G_i_j => 
                           C_6_port);
   G_L2_2_16_28 : g_block_2 port map( G_i_k => Gmat_28_17_port, G_kmin1_j => 
                           C_4_port, P_i_k => Pmat_28_17_port, G_i_j => 
                           C_7_port);
   G_L2_2_16_32 : g_block_1 port map( G_i_k => Gmat_32_17_port, G_kmin1_j => 
                           C_4_port, P_i_k => Pmat_32_17_port, G_i_j => 
                           C_8_port);
   U1 : INV_X1 port map( A => n2, ZN => n1);
   U2 : AOI21_X1 port map( B1 => P(0), B2 => Cin, A => G(0), ZN => n2);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity pg_network_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  P, G : out std_logic_vector
         (31 downto 0));

end pg_network_N32;

architecture SYN_ARCHDATAFLOW of pg_network_N32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B(9), B => A(9), Z => P(9));
   U2 : XOR2_X1 port map( A => B(8), B => A(8), Z => P(8));
   U3 : XOR2_X1 port map( A => B(7), B => A(7), Z => P(7));
   U4 : XOR2_X1 port map( A => B(6), B => A(6), Z => P(6));
   U5 : XOR2_X1 port map( A => B(5), B => A(5), Z => P(5));
   U6 : XOR2_X1 port map( A => B(4), B => A(4), Z => P(4));
   U7 : XOR2_X1 port map( A => B(3), B => A(3), Z => P(3));
   U8 : XOR2_X1 port map( A => B(31), B => A(31), Z => P(31));
   U9 : XOR2_X1 port map( A => B(30), B => A(30), Z => P(30));
   U10 : XOR2_X1 port map( A => B(2), B => A(2), Z => P(2));
   U11 : XOR2_X1 port map( A => B(29), B => A(29), Z => P(29));
   U12 : XOR2_X1 port map( A => B(28), B => A(28), Z => P(28));
   U13 : XOR2_X1 port map( A => B(27), B => A(27), Z => P(27));
   U14 : XOR2_X1 port map( A => B(26), B => A(26), Z => P(26));
   U15 : XOR2_X1 port map( A => B(25), B => A(25), Z => P(25));
   U16 : XOR2_X1 port map( A => B(24), B => A(24), Z => P(24));
   U17 : XOR2_X1 port map( A => B(23), B => A(23), Z => P(23));
   U18 : XOR2_X1 port map( A => B(22), B => A(22), Z => P(22));
   U19 : XOR2_X1 port map( A => B(21), B => A(21), Z => P(21));
   U20 : XOR2_X1 port map( A => B(20), B => A(20), Z => P(20));
   U21 : XOR2_X1 port map( A => B(1), B => A(1), Z => P(1));
   U22 : XOR2_X1 port map( A => B(19), B => A(19), Z => P(19));
   U23 : XOR2_X1 port map( A => B(18), B => A(18), Z => P(18));
   U24 : XOR2_X1 port map( A => B(17), B => A(17), Z => P(17));
   U25 : XOR2_X1 port map( A => B(16), B => A(16), Z => P(16));
   U26 : XOR2_X1 port map( A => B(15), B => A(15), Z => P(15));
   U27 : XOR2_X1 port map( A => B(14), B => A(14), Z => P(14));
   U28 : XOR2_X1 port map( A => B(13), B => A(13), Z => P(13));
   U29 : XOR2_X1 port map( A => B(12), B => A(12), Z => P(12));
   U30 : XOR2_X1 port map( A => B(11), B => A(11), Z => P(11));
   U31 : XOR2_X1 port map( A => B(10), B => A(10), Z => P(10));
   U32 : XOR2_X1 port map( A => B(0), B => A(0), Z => P(0));
   U33 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => G(9));
   U34 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => G(8));
   U35 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => G(7));
   U36 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => G(6));
   U37 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => G(5));
   U38 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => G(4));
   U39 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => G(3));
   U40 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => G(31));
   U41 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => G(30));
   U42 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => G(2));
   U43 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => G(29));
   U44 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => G(28));
   U45 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => G(27));
   U46 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => G(26));
   U47 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => G(25));
   U48 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => G(24));
   U49 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => G(23));
   U50 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => G(22));
   U51 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => G(21));
   U52 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => G(20));
   U53 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => G(1));
   U54 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => G(19));
   U55 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => G(18));
   U56 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => G(17));
   U57 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => G(16));
   U58 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => G(15));
   U59 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => G(14));
   U60 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => G(13));
   U61 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => G(12));
   U62 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => G(11));
   U63 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => G(10));
   U64 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => G(0));

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity sum_generator_N32_Nbit_blocks4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Carry 
         : in std_logic_vector (7 downto 0);  S : out std_logic_vector (31 
         downto 0);  Cout : out std_logic);

end sum_generator_N32_Nbit_blocks4;

architecture SYN_ARCHSTRUCT of sum_generator_N32_Nbit_blocks4 is

   component carry_select_block_N4_1
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_2
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_3
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_4
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_5
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_6
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_7
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_0
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   Cout <= Carry(7);
   
   CSB_1 : carry_select_block_N4_0 port map( Cin => Cin, A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(3) => B(3), B(2)
                           => B(2), B(1) => B(1), B(0) => B(0), S(3) => S(3), 
                           S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSB_2 : carry_select_block_N4_7 port map( Cin => Carry(0), A(3) => A(7), 
                           A(2) => A(6), A(1) => A(5), A(0) => A(4), B(3) => 
                           B(7), B(2) => B(6), B(1) => B(5), B(0) => B(4), S(3)
                           => S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CSB_3 : carry_select_block_N4_6 port map( Cin => Carry(1), A(3) => A(11), 
                           A(2) => A(10), A(1) => A(9), A(0) => A(8), B(3) => 
                           B(11), B(2) => B(10), B(1) => B(9), B(0) => B(8), 
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   CSB_4 : carry_select_block_N4_5 port map( Cin => Carry(2), A(3) => A(15), 
                           A(2) => A(14), A(1) => A(13), A(0) => A(12), B(3) =>
                           B(15), B(2) => B(14), B(1) => B(13), B(0) => B(12), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));
   CSB_5 : carry_select_block_N4_4 port map( Cin => Carry(3), A(3) => A(19), 
                           A(2) => A(18), A(1) => A(17), A(0) => A(16), B(3) =>
                           B(19), B(2) => B(18), B(1) => B(17), B(0) => B(16), 
                           S(3) => S(19), S(2) => S(18), S(1) => S(17), S(0) =>
                           S(16));
   CSB_6 : carry_select_block_N4_3 port map( Cin => Carry(4), A(3) => A(23), 
                           A(2) => A(22), A(1) => A(21), A(0) => A(20), B(3) =>
                           B(23), B(2) => B(22), B(1) => B(21), B(0) => B(20), 
                           S(3) => S(23), S(2) => S(22), S(1) => S(21), S(0) =>
                           S(20));
   CSB_7 : carry_select_block_N4_2 port map( Cin => Carry(5), A(3) => A(27), 
                           A(2) => A(26), A(1) => A(25), A(0) => A(24), B(3) =>
                           B(27), B(2) => B(26), B(1) => B(25), B(0) => B(24), 
                           S(3) => S(27), S(2) => S(26), S(1) => S(25), S(0) =>
                           S(24));
   CSB_8 : carry_select_block_N4_1 port map( Cin => Carry(6), A(3) => A(31), 
                           A(2) => A(30), A(1) => A(29), A(0) => A(28), B(3) =>
                           B(31), B(2) => B(30), B(1) => B(29), B(0) => B(28), 
                           S(3) => S(31), S(2) => S(30), S(1) => S(29), S(0) =>
                           S(28));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity carry_generator_N32_carry_range4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  C : 
         out std_logic_vector (8 downto 0));

end carry_generator_N32_carry_range4;

architecture SYN_ARCHSTRUCT of carry_generator_N32_carry_range4 is

   component carry_generator_sparse_tree_N32_carry_range4
      port( P, G : in std_logic_vector (31 downto 0);  Cin : in std_logic;  C :
            out std_logic_vector (8 downto 0));
   end component;
   
   component pg_network_N32
      port( A, B : in std_logic_vector (31 downto 0);  P, G : out 
            std_logic_vector (31 downto 0));
   end component;
   
   signal P_31_port, P_30_port, P_29_port, P_28_port, P_27_port, P_26_port, 
      P_25_port, P_24_port, P_23_port, P_22_port, P_21_port, P_20_port, 
      P_19_port, P_18_port, P_17_port, P_16_port, P_15_port, P_14_port, 
      P_13_port, P_12_port, P_11_port, P_10_port, P_9_port, P_8_port, P_7_port,
      P_6_port, P_5_port, P_4_port, P_3_port, P_2_port, P_1_port, P_0_port, 
      G_31_port, G_30_port, G_29_port, G_28_port, G_27_port, G_26_port, 
      G_25_port, G_24_port, G_23_port, G_22_port, G_21_port, G_20_port, 
      G_19_port, G_18_port, G_17_port, G_16_port, G_15_port, G_14_port, 
      G_13_port, G_12_port, G_11_port, G_10_port, G_9_port, G_8_port, G_7_port,
      G_6_port, G_5_port, G_4_port, G_3_port, G_2_port, G_1_port, G_0_port : 
      std_logic;

begin
   
   PG_NET : pg_network_N32 port map( A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), P(31) => P_31_port, P(30) => P_30_port, 
                           P(29) => P_29_port, P(28) => P_28_port, P(27) => 
                           P_27_port, P(26) => P_26_port, P(25) => P_25_port, 
                           P(24) => P_24_port, P(23) => P_23_port, P(22) => 
                           P_22_port, P(21) => P_21_port, P(20) => P_20_port, 
                           P(19) => P_19_port, P(18) => P_18_port, P(17) => 
                           P_17_port, P(16) => P_16_port, P(15) => P_15_port, 
                           P(14) => P_14_port, P(13) => P_13_port, P(12) => 
                           P_12_port, P(11) => P_11_port, P(10) => P_10_port, 
                           P(9) => P_9_port, P(8) => P_8_port, P(7) => P_7_port
                           , P(6) => P_6_port, P(5) => P_5_port, P(4) => 
                           P_4_port, P(3) => P_3_port, P(2) => P_2_port, P(1) 
                           => P_1_port, P(0) => P_0_port, G(31) => G_31_port, 
                           G(30) => G_30_port, G(29) => G_29_port, G(28) => 
                           G_28_port, G(27) => G_27_port, G(26) => G_26_port, 
                           G(25) => G_25_port, G(24) => G_24_port, G(23) => 
                           G_23_port, G(22) => G_22_port, G(21) => G_21_port, 
                           G(20) => G_20_port, G(19) => G_19_port, G(18) => 
                           G_18_port, G(17) => G_17_port, G(16) => G_16_port, 
                           G(15) => G_15_port, G(14) => G_14_port, G(13) => 
                           G_13_port, G(12) => G_12_port, G(11) => G_11_port, 
                           G(10) => G_10_port, G(9) => G_9_port, G(8) => 
                           G_8_port, G(7) => G_7_port, G(6) => G_6_port, G(5) 
                           => G_5_port, G(4) => G_4_port, G(3) => G_3_port, 
                           G(2) => G_2_port, G(1) => G_1_port, G(0) => G_0_port
                           );
   CG : carry_generator_sparse_tree_N32_carry_range4 port map( P(31) => 
                           P_31_port, P(30) => P_30_port, P(29) => P_29_port, 
                           P(28) => P_28_port, P(27) => P_27_port, P(26) => 
                           P_26_port, P(25) => P_25_port, P(24) => P_24_port, 
                           P(23) => P_23_port, P(22) => P_22_port, P(21) => 
                           P_21_port, P(20) => P_20_port, P(19) => P_19_port, 
                           P(18) => P_18_port, P(17) => P_17_port, P(16) => 
                           P_16_port, P(15) => P_15_port, P(14) => P_14_port, 
                           P(13) => P_13_port, P(12) => P_12_port, P(11) => 
                           P_11_port, P(10) => P_10_port, P(9) => P_9_port, 
                           P(8) => P_8_port, P(7) => P_7_port, P(6) => P_6_port
                           , P(5) => P_5_port, P(4) => P_4_port, P(3) => 
                           P_3_port, P(2) => P_2_port, P(1) => P_1_port, P(0) 
                           => P_0_port, G(31) => G_31_port, G(30) => G_30_port,
                           G(29) => G_29_port, G(28) => G_28_port, G(27) => 
                           G_27_port, G(26) => G_26_port, G(25) => G_25_port, 
                           G(24) => G_24_port, G(23) => G_23_port, G(22) => 
                           G_22_port, G(21) => G_21_port, G(20) => G_20_port, 
                           G(19) => G_19_port, G(18) => G_18_port, G(17) => 
                           G_17_port, G(16) => G_16_port, G(15) => G_15_port, 
                           G(14) => G_14_port, G(13) => G_13_port, G(12) => 
                           G_12_port, G(11) => G_11_port, G(10) => G_10_port, 
                           G(9) => G_9_port, G(8) => G_8_port, G(7) => G_7_port
                           , G(6) => G_6_port, G(5) => G_5_port, G(4) => 
                           G_4_port, G(3) => G_3_port, G(2) => G_2_port, G(1) 
                           => G_1_port, G(0) => G_0_port, Cin => Cin, C(8) => 
                           C(8), C(7) => C(7), C(6) => C(6), C(5) => C(5), C(4)
                           => C(4), C(3) => C(3), C(2) => C(2), C(1) => C(1), 
                           C(0) => C(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_P4_adder_Nbit_blocks4.all;

entity P4_adder_Nbit_blocks4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4_adder_Nbit_blocks4;

architecture SYN_STRUCT of P4_adder_Nbit_blocks4 is

   component sum_generator_N32_Nbit_blocks4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  
            Carry : in std_logic_vector (7 downto 0);  S : out std_logic_vector
            (31 downto 0);  Cout : out std_logic);
   end component;
   
   component carry_generator_N32_carry_range4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  C :
            out std_logic_vector (8 downto 0));
   end component;
   
   signal Carries_8_port, Carries_7_port, Carries_6_port, Carries_5_port, 
      Carries_4_port, Carries_3_port, Carries_2_port, Carries_1_port, n_1016 : 
      std_logic;

begin
   
   CG : carry_generator_N32_carry_range4 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Cin => Cin, C(8) => 
                           Carries_8_port, C(7) => Carries_7_port, C(6) => 
                           Carries_6_port, C(5) => Carries_5_port, C(4) => 
                           Carries_4_port, C(3) => Carries_3_port, C(2) => 
                           Carries_2_port, C(1) => Carries_1_port, C(0) => 
                           n_1016);
   SG : sum_generator_N32_Nbit_blocks4 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Cin => Cin, Carry(7) => 
                           Carries_8_port, Carry(6) => Carries_7_port, Carry(5)
                           => Carries_6_port, Carry(4) => Carries_5_port, 
                           Carry(3) => Carries_4_port, Carry(2) => 
                           Carries_3_port, Carry(1) => Carries_2_port, Carry(0)
                           => Carries_1_port, S(31) => S(31), S(30) => S(30), 
                           S(29) => S(29), S(28) => S(28), S(27) => S(27), 
                           S(26) => S(26), S(25) => S(25), S(24) => S(24), 
                           S(23) => S(23), S(22) => S(22), S(21) => S(21), 
                           S(20) => S(20), S(19) => S(19), S(18) => S(18), 
                           S(17) => S(17), S(16) => S(16), S(15) => S(15), 
                           S(14) => S(14), S(13) => S(13), S(12) => S(12), 
                           S(11) => S(11), S(10) => S(10), S(9) => S(9), S(8) 
                           => S(8), S(7) => S(7), S(6) => S(6), S(5) => S(5), 
                           S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1) => 
                           S(1), S(0) => S(0), Cout => Cout);

end SYN_STRUCT;
