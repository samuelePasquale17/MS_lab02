library ieee;
use ieee.std_logic_1164.all;
use work.constants.all;

entity carry_select_block is
    generic (
        N : integer := Nbit_carry_select_block     -- size Number of Bits
    );
    port (
        Cin : in std_logic;
        A : in std_logic_vector(N-1 downto 0);
        B : in std_logic_vector(N-1 downto 0);
        S : out std_logic_vector(N-1 downto 0)
    );
end carry_select_block;

architecture ARCHSTRUCT of carry_select_block is

    -- RCA component
    component RCA is
        generic (
            DRCAS 	: time 		:= DelaySum_RCA;		
            DRCAC 	: time 		:= DelayCarryOut_RCA;		
            N 	: integer 	    := Nbit_carry_select_block
        );
        port(
            A 	: 	in 		std_logic_vector(N-1 downto 0);
            B 	: 	in 		std_logic_vector(N-1 downto 0);
            Ci 	: 	in 		std_logic;
            S 	: 	out 	std_logic_vector(N-1 downto 0);
            Co 	: 	out 	std_logic
        );
    end component;

    component muxN1 is
        generic (
            N : integer := Nbit_carry_select_block
        );
        port (
			A : 	in 		std_logic_vector(N-1 downto 0);
			B : 	in 		std_logic_vector(N-1 downto 0);
			S : 	in 		std_logic;
			Y : 	out 	std_logic_vector(N-1 downto 0)
        );
    end component;

    signal S1, S2 : std_logic_vector(N-1 downto 0); -- sum generated by RCAs

begin

    -- RCA n.1 with Carry In set to 0
    RCA1 : RCA 
    generic map(DRCAS => DelaySum_RCA, DRCAC => DelayCarryOut_RCA, N => Nbit_carry_select_block)
    port map(A => A, B => B, Ci => '0', S => S1, Co => open);

    -- RCA n.2 with Carry In set to 1
    RCA2 : RCA 
    generic map(DRCAS => DelaySum_RCA, DRCAC => DelayCarryOut_RCA, N => Nbit_carry_select_block)
    port map(A => A, B => B, Ci => '1', S => S2, Co => open);

    MUX : muxN1
    generic map(N => N)       -- if carry in is '0' B is driven as output,
    port map(A => S2, B => S1, S => Cin, Y => S);   -- otherwise A is the MUX outcome 

end architecture;

configuration CFG_CARRY_SELECT_BLOCK_ARCHSTRUCT of carry_select_block is
    for ARCHSTRUCT
        for all : RCA 
            use configuration work.CFG_RCA_ARCHSTRUCT;
        end for;

        for MUX : muxN1 
            use configuration work.CFG_MUXN1_ARCHSTRUCT;
        end for;
    end for;

end configuration;
