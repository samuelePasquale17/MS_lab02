
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL_N8 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL_N8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_0_DW01_add_0_DW01_add_7 is

   port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (13 downto 0);  CO : out std_logic);

end shift_pow2_N8_0_DW01_add_0_DW01_add_7;

architecture SYN_cla of shift_pow2_N8_0_DW01_add_0_DW01_add_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, n1, SUM_7_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SUM <= ( SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, SUM_7_port, A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n1);
   U3 : INV_X1 port map( A => n12, ZN => n7);
   U4 : INV_X1 port map( A => n24, ZN => n4);
   U5 : INV_X1 port map( A => n27, ZN => n5);
   U6 : INV_X1 port map( A => n16, ZN => n8);
   U7 : INV_X1 port map( A => n32, ZN => n6);
   U8 : INV_X1 port map( A => n20, ZN => n3);
   U9 : XNOR2_X1 port map( A => B(13), B => n17, ZN => SUM_13_port);
   U10 : AND2_X1 port map( A1 => n16, A2 => n1, ZN => SUM_7_port);
   U11 : XNOR2_X1 port map( A => n9, B => n10, ZN => SUM_9_port);
   U12 : NOR2_X1 port map( A1 => n7, A2 => n11, ZN => n10);
   U13 : XOR2_X1 port map( A => n8, B => n13, Z => SUM_8_port);
   U14 : AND2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U15 : AOI21_X1 port map( B1 => n18, B2 => n3, A => n19, ZN => n17);
   U16 : XOR2_X1 port map( A => n18, B => n21, Z => SUM_12_port);
   U17 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U18 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n19);
   U19 : NOR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n20);
   U20 : OAI211_X1 port map( C1 => n22, C2 => n23, A => n24, B => n25, ZN => 
                           n18);
   U21 : OR4_X1 port map( A1 => n26, A2 => n27, A3 => n23, A4 => n11, ZN => n25
                           );
   U22 : AOI21_X1 port map( B1 => n5, B2 => n28, A => n6, ZN => n22);
   U23 : OAI21_X1 port map( B1 => n11, B2 => n15, A => n12, ZN => n28);
   U24 : XNOR2_X1 port map( A => n29, B => n30, ZN => SUM_11_port);
   U25 : NOR2_X1 port map( A1 => n23, A2 => n4, ZN => n30);
   U26 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n24);
   U27 : NOR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n23);
   U28 : AOI21_X1 port map( B1 => n31, B2 => n5, A => n6, ZN => n29);
   U29 : XNOR2_X1 port map( A => n33, B => n31, ZN => SUM_10_port);
   U30 : OAI21_X1 port map( B1 => n11, B2 => n9, A => n12, ZN => n31);
   U31 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n12);
   U32 : AND2_X1 port map( A1 => n26, A2 => n15, ZN => n9);
   U33 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n15);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n14, ZN => n26);
   U35 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n14);
   U36 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n16);
   U37 : NOR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n11);
   U38 : NAND2_X1 port map( A1 => n32, A2 => n5, ZN => n33);
   U39 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n27);
   U40 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n32);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_0_DW02_mult_0_DW02_mult_7 is

   port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  PRODUCT 
         : out std_logic_vector (15 downto 0));

end shift_pow2_N8_0_DW02_mult_0_DW02_mult_7;

architecture SYN_csa of shift_pow2_N8_0_DW02_mult_0_DW02_mult_7 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component shift_pow2_N8_0_DW01_add_0_DW01_add_7
      port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (13 downto 0);  CO : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, ab_7_4_port, 
      ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_7_port, ab_3_6_port, 
      ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, 
      ab_3_0_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, ab_2_4_port, 
      ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, ab_1_7_port, 
      ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_2_port, 
      ab_1_1_port, ab_1_0_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, 
      SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, SUMB_7_0_port, SUMB_6_6_port
      , SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, 
      SUMB_6_1_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_6_port, SUMB_4_5_port, 
      SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_6_port
      , SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, 
      SUMB_3_1_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n_1011 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => 
                           SUMB_7_0_port);
   S4_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S4_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S4_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S4_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S4_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S5_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           ab_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S3_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           ab_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S3_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           ab_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S3_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           ab_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S3_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           ab_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n7, CI => n14, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n6, CI => n13, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n5, CI => n12, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n4, CI => n11, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n3, CI => n10, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n2, CI => n9, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S3_2_6 : FA_X1 port map( A => ab_2_6_port, B => n8, CI => ab_1_7_port, CO =>
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   FS_1 : shift_pow2_N8_0_DW01_add_0_DW01_add_7 port map( A(13) => n46, A(12) 
                           => n18, A(11) => n21, A(10) => n19, A(9) => n22, 
                           A(8) => n27, A(7) => n20, A(6) => n17, A(5) => 
                           SUMB_7_0_port, A(4) => A1_4_port, A(3) => A1_3_port,
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(13) => n15, B(12) => n28, B(11) => n25,
                           B(10) => n24, B(9) => n26, B(8) => n29, B(7) => n23,
                           B(6) => n46, B(5) => n47, B(4) => n47, B(3) => n47, 
                           B(2) => n47, B(1) => n47, B(0) => X_Logic0_port, CI 
                           => X_Logic0_port, SUM(13) => PRODUCT(15), SUM(12) =>
                           PRODUCT(14), SUM(11) => PRODUCT(13), SUM(10) => 
                           PRODUCT(12), SUM(9) => PRODUCT(11), SUM(8) => 
                           PRODUCT(10), SUM(7) => PRODUCT(9), SUM(6) => 
                           PRODUCT(8), SUM(5) => PRODUCT(7), SUM(4) => 
                           PRODUCT(6), SUM(3) => PRODUCT(5), SUM(2) => 
                           PRODUCT(4), SUM(1) => PRODUCT(3), SUM(0) => 
                           PRODUCT(2), CO => n_1011);
   U2 : INV_X1 port map( A => B(4), ZN => n35);
   U3 : INV_X1 port map( A => B(5), ZN => n34);
   U4 : INV_X1 port map( A => B(6), ZN => n33);
   U5 : INV_X1 port map( A => B(7), ZN => n30);
   U6 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n2);
   U7 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n3);
   U8 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n4);
   U9 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n5);
   U10 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n6);
   U11 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n7);
   U12 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n8);
   U13 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n9);
   U14 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n10);
   U15 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n11);
   U16 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n12);
   U17 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n13);
   U18 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n14);
   U19 : AND2_X1 port map( A1 => CARRYB_7_6_port, A2 => ab_7_7_port, ZN => n15)
                           ;
   U20 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U21 : XOR2_X1 port map( A => CARRYB_7_0_port, B => SUMB_7_1_port, Z => n17);
   U22 : XOR2_X1 port map( A => CARRYB_7_6_port, B => ab_7_7_port, Z => n18);
   U23 : XOR2_X1 port map( A => CARRYB_7_4_port, B => SUMB_7_5_port, Z => n19);
   U24 : XOR2_X1 port map( A => CARRYB_7_1_port, B => SUMB_7_2_port, Z => n20);
   U25 : XOR2_X1 port map( A => CARRYB_7_5_port, B => SUMB_7_6_port, Z => n21);
   U26 : XOR2_X1 port map( A => CARRYB_7_3_port, B => SUMB_7_4_port, Z => n22);
   U27 : AND2_X1 port map( A1 => CARRYB_7_0_port, A2 => SUMB_7_1_port, ZN => 
                           n23);
   U28 : AND2_X1 port map( A1 => CARRYB_7_3_port, A2 => SUMB_7_4_port, ZN => 
                           n24);
   U29 : AND2_X1 port map( A1 => CARRYB_7_4_port, A2 => SUMB_7_5_port, ZN => 
                           n25);
   U30 : AND2_X1 port map( A1 => CARRYB_7_2_port, A2 => SUMB_7_3_port, ZN => 
                           n26);
   U31 : XOR2_X1 port map( A => CARRYB_7_2_port, B => SUMB_7_3_port, Z => n27);
   U32 : AND2_X1 port map( A1 => CARRYB_7_5_port, A2 => SUMB_7_6_port, ZN => 
                           n28);
   U33 : AND2_X1 port map( A1 => CARRYB_7_1_port, A2 => SUMB_7_2_port, ZN => 
                           n29);
   U34 : INV_X1 port map( A => B(3), ZN => n31);
   U35 : INV_X1 port map( A => B(2), ZN => n32);
   U36 : INV_X1 port map( A => B(1), ZN => n36);
   U37 : INV_X1 port map( A => B(0), ZN => n37);
   U38 : INV_X1 port map( A => A(7), ZN => n38);
   U39 : INV_X1 port map( A => A(0), ZN => n45);
   U40 : INV_X1 port map( A => A(1), ZN => n44);
   U41 : INV_X1 port map( A => A(3), ZN => n42);
   U42 : INV_X1 port map( A => A(4), ZN => n41);
   U43 : INV_X1 port map( A => A(5), ZN => n40);
   U44 : INV_X1 port map( A => A(6), ZN => n39);
   U45 : INV_X1 port map( A => A(2), ZN => n43);
   n46 <= '0';
   U47 : NOR2_X1 port map( A1 => n38, A2 => n30, ZN => ab_7_7_port);
   U48 : NOR2_X1 port map( A1 => n38, A2 => n33, ZN => ab_7_6_port);
   U49 : NOR2_X1 port map( A1 => n38, A2 => n34, ZN => ab_7_5_port);
   U50 : NOR2_X1 port map( A1 => n38, A2 => n35, ZN => ab_7_4_port);
   U51 : NOR2_X1 port map( A1 => n38, A2 => n31, ZN => ab_7_3_port);
   U52 : NOR2_X1 port map( A1 => n38, A2 => n32, ZN => ab_7_2_port);
   U53 : NOR2_X1 port map( A1 => n38, A2 => n36, ZN => ab_7_1_port);
   U54 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => ab_7_0_port);
   U55 : NOR2_X1 port map( A1 => n30, A2 => n39, ZN => ab_6_7_port);
   U56 : NOR2_X1 port map( A1 => n33, A2 => n39, ZN => ab_6_6_port);
   U57 : NOR2_X1 port map( A1 => n34, A2 => n39, ZN => ab_6_5_port);
   U58 : NOR2_X1 port map( A1 => n35, A2 => n39, ZN => ab_6_4_port);
   U59 : NOR2_X1 port map( A1 => n31, A2 => n39, ZN => ab_6_3_port);
   U60 : NOR2_X1 port map( A1 => n32, A2 => n39, ZN => ab_6_2_port);
   U61 : NOR2_X1 port map( A1 => n36, A2 => n39, ZN => ab_6_1_port);
   U62 : NOR2_X1 port map( A1 => n37, A2 => n39, ZN => ab_6_0_port);
   U63 : NOR2_X1 port map( A1 => n30, A2 => n40, ZN => ab_5_7_port);
   U64 : NOR2_X1 port map( A1 => n33, A2 => n40, ZN => ab_5_6_port);
   U65 : NOR2_X1 port map( A1 => n34, A2 => n40, ZN => ab_5_5_port);
   U66 : NOR2_X1 port map( A1 => n35, A2 => n40, ZN => ab_5_4_port);
   U67 : NOR2_X1 port map( A1 => n31, A2 => n40, ZN => ab_5_3_port);
   U68 : NOR2_X1 port map( A1 => n32, A2 => n40, ZN => ab_5_2_port);
   U69 : NOR2_X1 port map( A1 => n36, A2 => n40, ZN => ab_5_1_port);
   U70 : NOR2_X1 port map( A1 => n37, A2 => n40, ZN => ab_5_0_port);
   U71 : NOR2_X1 port map( A1 => n30, A2 => n41, ZN => ab_4_7_port);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n41, ZN => ab_4_6_port);
   U73 : NOR2_X1 port map( A1 => n34, A2 => n41, ZN => ab_4_5_port);
   U74 : NOR2_X1 port map( A1 => n35, A2 => n41, ZN => ab_4_4_port);
   U75 : NOR2_X1 port map( A1 => n31, A2 => n41, ZN => ab_4_3_port);
   U76 : NOR2_X1 port map( A1 => n32, A2 => n41, ZN => ab_4_2_port);
   U77 : NOR2_X1 port map( A1 => n36, A2 => n41, ZN => ab_4_1_port);
   U78 : NOR2_X1 port map( A1 => n37, A2 => n41, ZN => ab_4_0_port);
   U79 : NOR2_X1 port map( A1 => n30, A2 => n42, ZN => ab_3_7_port);
   U80 : NOR2_X1 port map( A1 => n33, A2 => n42, ZN => ab_3_6_port);
   U81 : NOR2_X1 port map( A1 => n34, A2 => n42, ZN => ab_3_5_port);
   U82 : NOR2_X1 port map( A1 => n35, A2 => n42, ZN => ab_3_4_port);
   U83 : NOR2_X1 port map( A1 => n31, A2 => n42, ZN => ab_3_3_port);
   U84 : NOR2_X1 port map( A1 => n32, A2 => n42, ZN => ab_3_2_port);
   U85 : NOR2_X1 port map( A1 => n36, A2 => n42, ZN => ab_3_1_port);
   U86 : NOR2_X1 port map( A1 => n37, A2 => n42, ZN => ab_3_0_port);
   U87 : NOR2_X1 port map( A1 => n30, A2 => n43, ZN => ab_2_7_port);
   U88 : NOR2_X1 port map( A1 => n33, A2 => n43, ZN => ab_2_6_port);
   U89 : NOR2_X1 port map( A1 => n34, A2 => n43, ZN => ab_2_5_port);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n43, ZN => ab_2_4_port);
   U91 : NOR2_X1 port map( A1 => n31, A2 => n43, ZN => ab_2_3_port);
   U92 : NOR2_X1 port map( A1 => n32, A2 => n43, ZN => ab_2_2_port);
   U93 : NOR2_X1 port map( A1 => n36, A2 => n43, ZN => ab_2_1_port);
   U94 : NOR2_X1 port map( A1 => n37, A2 => n43, ZN => ab_2_0_port);
   U95 : NOR2_X1 port map( A1 => n30, A2 => n44, ZN => ab_1_7_port);
   U96 : NOR2_X1 port map( A1 => n33, A2 => n44, ZN => ab_1_6_port);
   U97 : NOR2_X1 port map( A1 => n34, A2 => n44, ZN => ab_1_5_port);
   U98 : NOR2_X1 port map( A1 => n35, A2 => n44, ZN => ab_1_4_port);
   U99 : NOR2_X1 port map( A1 => n31, A2 => n44, ZN => ab_1_3_port);
   U100 : NOR2_X1 port map( A1 => n32, A2 => n44, ZN => ab_1_2_port);
   U101 : NOR2_X1 port map( A1 => n36, A2 => n44, ZN => ab_1_1_port);
   U102 : NOR2_X1 port map( A1 => n37, A2 => n44, ZN => ab_1_0_port);
   U103 : NOR2_X1 port map( A1 => n30, A2 => n45, ZN => ab_0_7_port);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n45, ZN => ab_0_6_port);
   U105 : NOR2_X1 port map( A1 => n34, A2 => n45, ZN => ab_0_5_port);
   U106 : NOR2_X1 port map( A1 => n35, A2 => n45, ZN => ab_0_4_port);
   U107 : NOR2_X1 port map( A1 => n31, A2 => n45, ZN => ab_0_3_port);
   U108 : NOR2_X1 port map( A1 => n32, A2 => n45, ZN => ab_0_2_port);
   U109 : NOR2_X1 port map( A1 => n36, A2 => n45, ZN => ab_0_1_port);
   U110 : NOR2_X1 port map( A1 => n37, A2 => n45, ZN => PRODUCT(0));
   n47 <= '0';

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_7_DW01_add_0_DW01_add_6 is

   port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (13 downto 0);  CO : out std_logic);

end shift_pow2_N8_7_DW01_add_0_DW01_add_6;

architecture SYN_cla of shift_pow2_N8_7_DW01_add_0_DW01_add_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, n1, SUM_7_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SUM <= ( SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, SUM_7_port, A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n1);
   U3 : INV_X1 port map( A => n12, ZN => n7);
   U4 : INV_X1 port map( A => n24, ZN => n4);
   U5 : INV_X1 port map( A => n27, ZN => n5);
   U6 : INV_X1 port map( A => n16, ZN => n8);
   U7 : INV_X1 port map( A => n32, ZN => n6);
   U8 : INV_X1 port map( A => n20, ZN => n3);
   U9 : XNOR2_X1 port map( A => B(13), B => n17, ZN => SUM_13_port);
   U10 : AND2_X1 port map( A1 => n16, A2 => n1, ZN => SUM_7_port);
   U11 : XNOR2_X1 port map( A => n9, B => n10, ZN => SUM_9_port);
   U12 : NOR2_X1 port map( A1 => n7, A2 => n11, ZN => n10);
   U13 : XOR2_X1 port map( A => n8, B => n13, Z => SUM_8_port);
   U14 : AND2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U15 : AOI21_X1 port map( B1 => n18, B2 => n3, A => n19, ZN => n17);
   U16 : XOR2_X1 port map( A => n18, B => n21, Z => SUM_12_port);
   U17 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U18 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n19);
   U19 : NOR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n20);
   U20 : OAI211_X1 port map( C1 => n22, C2 => n23, A => n24, B => n25, ZN => 
                           n18);
   U21 : OR4_X1 port map( A1 => n26, A2 => n27, A3 => n23, A4 => n11, ZN => n25
                           );
   U22 : AOI21_X1 port map( B1 => n5, B2 => n28, A => n6, ZN => n22);
   U23 : OAI21_X1 port map( B1 => n11, B2 => n15, A => n12, ZN => n28);
   U24 : XNOR2_X1 port map( A => n29, B => n30, ZN => SUM_11_port);
   U25 : NOR2_X1 port map( A1 => n23, A2 => n4, ZN => n30);
   U26 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n24);
   U27 : NOR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n23);
   U28 : AOI21_X1 port map( B1 => n31, B2 => n5, A => n6, ZN => n29);
   U29 : XNOR2_X1 port map( A => n33, B => n31, ZN => SUM_10_port);
   U30 : OAI21_X1 port map( B1 => n11, B2 => n9, A => n12, ZN => n31);
   U31 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n12);
   U32 : AND2_X1 port map( A1 => n26, A2 => n15, ZN => n9);
   U33 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n15);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n14, ZN => n26);
   U35 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n14);
   U36 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n16);
   U37 : NOR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n11);
   U38 : NAND2_X1 port map( A1 => n32, A2 => n5, ZN => n33);
   U39 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n27);
   U40 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n32);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_7_DW02_mult_0_DW02_mult_6 is

   port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  PRODUCT 
         : out std_logic_vector (15 downto 0));

end shift_pow2_N8_7_DW02_mult_0_DW02_mult_6;

architecture SYN_csa of shift_pow2_N8_7_DW02_mult_0_DW02_mult_6 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component shift_pow2_N8_7_DW01_add_0_DW01_add_6
      port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (13 downto 0);  CO : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, ab_7_4_port, 
      ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_7_port, ab_3_6_port, 
      ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, 
      ab_3_0_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, ab_2_4_port, 
      ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, ab_1_7_port, 
      ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_2_port, 
      ab_1_1_port, ab_1_0_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, 
      SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, SUMB_7_0_port, SUMB_6_6_port
      , SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, 
      SUMB_6_1_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_6_port, SUMB_4_5_port, 
      SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_6_port
      , SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, 
      SUMB_3_1_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n_1023 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => 
                           SUMB_7_0_port);
   S4_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S4_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S4_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S4_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S4_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S5_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           ab_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S3_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           ab_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S3_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           ab_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S3_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           ab_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S3_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           ab_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n7, CI => n14, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n6, CI => n13, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n5, CI => n12, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n4, CI => n11, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n3, CI => n10, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n2, CI => n9, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S3_2_6 : FA_X1 port map( A => ab_2_6_port, B => n8, CI => ab_1_7_port, CO =>
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   FS_1 : shift_pow2_N8_7_DW01_add_0_DW01_add_6 port map( A(13) => n46, A(12) 
                           => n17, A(11) => n21, A(10) => n19, A(9) => n22, 
                           A(8) => n27, A(7) => n20, A(6) => n18, A(5) => 
                           SUMB_7_0_port, A(4) => A1_4_port, A(3) => A1_3_port,
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(13) => n15, B(12) => n29, B(11) => n25,
                           B(10) => n24, B(9) => n26, B(8) => n28, B(7) => n23,
                           B(6) => n46, B(5) => n47, B(4) => n47, B(3) => n47, 
                           B(2) => n47, B(1) => n47, B(0) => X_Logic0_port, CI 
                           => X_Logic0_port, SUM(13) => PRODUCT(15), SUM(12) =>
                           PRODUCT(14), SUM(11) => PRODUCT(13), SUM(10) => 
                           PRODUCT(12), SUM(9) => PRODUCT(11), SUM(8) => 
                           PRODUCT(10), SUM(7) => PRODUCT(9), SUM(6) => 
                           PRODUCT(8), SUM(5) => PRODUCT(7), SUM(4) => 
                           PRODUCT(6), SUM(3) => PRODUCT(5), SUM(2) => 
                           PRODUCT(4), SUM(1) => PRODUCT(3), SUM(0) => 
                           PRODUCT(2), CO => n_1023);
   U2 : INV_X1 port map( A => B(4), ZN => n35);
   U3 : INV_X1 port map( A => B(5), ZN => n34);
   U4 : INV_X1 port map( A => B(6), ZN => n33);
   U5 : INV_X1 port map( A => B(7), ZN => n30);
   U6 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n2);
   U7 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n3);
   U8 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n4);
   U9 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n5);
   U10 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n6);
   U11 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n7);
   U12 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n8);
   U13 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n9);
   U14 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n10);
   U15 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n11);
   U16 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n12);
   U17 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n13);
   U18 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n14);
   U19 : AND2_X1 port map( A1 => CARRYB_7_6_port, A2 => ab_7_7_port, ZN => n15)
                           ;
   U20 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U21 : XOR2_X1 port map( A => CARRYB_7_6_port, B => ab_7_7_port, Z => n17);
   U22 : XOR2_X1 port map( A => CARRYB_7_0_port, B => SUMB_7_1_port, Z => n18);
   U23 : XOR2_X1 port map( A => CARRYB_7_4_port, B => SUMB_7_5_port, Z => n19);
   U24 : XOR2_X1 port map( A => CARRYB_7_1_port, B => SUMB_7_2_port, Z => n20);
   U25 : XOR2_X1 port map( A => CARRYB_7_5_port, B => SUMB_7_6_port, Z => n21);
   U26 : XOR2_X1 port map( A => CARRYB_7_3_port, B => SUMB_7_4_port, Z => n22);
   U27 : AND2_X1 port map( A1 => CARRYB_7_0_port, A2 => SUMB_7_1_port, ZN => 
                           n23);
   U28 : AND2_X1 port map( A1 => CARRYB_7_3_port, A2 => SUMB_7_4_port, ZN => 
                           n24);
   U29 : AND2_X1 port map( A1 => CARRYB_7_4_port, A2 => SUMB_7_5_port, ZN => 
                           n25);
   U30 : AND2_X1 port map( A1 => CARRYB_7_2_port, A2 => SUMB_7_3_port, ZN => 
                           n26);
   U31 : XOR2_X1 port map( A => CARRYB_7_2_port, B => SUMB_7_3_port, Z => n27);
   U32 : AND2_X1 port map( A1 => CARRYB_7_1_port, A2 => SUMB_7_2_port, ZN => 
                           n28);
   U33 : AND2_X1 port map( A1 => CARRYB_7_5_port, A2 => SUMB_7_6_port, ZN => 
                           n29);
   U34 : INV_X1 port map( A => B(3), ZN => n31);
   U35 : INV_X1 port map( A => B(2), ZN => n32);
   U36 : INV_X1 port map( A => B(1), ZN => n36);
   U37 : INV_X1 port map( A => B(0), ZN => n37);
   U38 : INV_X1 port map( A => A(7), ZN => n38);
   U39 : INV_X1 port map( A => A(0), ZN => n45);
   U40 : INV_X1 port map( A => A(1), ZN => n44);
   U41 : INV_X1 port map( A => A(3), ZN => n42);
   U42 : INV_X1 port map( A => A(2), ZN => n43);
   U43 : INV_X1 port map( A => A(4), ZN => n41);
   U44 : INV_X1 port map( A => A(5), ZN => n40);
   U45 : INV_X1 port map( A => A(6), ZN => n39);
   n46 <= '0';
   U47 : NOR2_X1 port map( A1 => n38, A2 => n30, ZN => ab_7_7_port);
   U48 : NOR2_X1 port map( A1 => n38, A2 => n33, ZN => ab_7_6_port);
   U49 : NOR2_X1 port map( A1 => n38, A2 => n34, ZN => ab_7_5_port);
   U50 : NOR2_X1 port map( A1 => n38, A2 => n35, ZN => ab_7_4_port);
   U51 : NOR2_X1 port map( A1 => n38, A2 => n31, ZN => ab_7_3_port);
   U52 : NOR2_X1 port map( A1 => n38, A2 => n32, ZN => ab_7_2_port);
   U53 : NOR2_X1 port map( A1 => n38, A2 => n36, ZN => ab_7_1_port);
   U54 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => ab_7_0_port);
   U55 : NOR2_X1 port map( A1 => n30, A2 => n39, ZN => ab_6_7_port);
   U56 : NOR2_X1 port map( A1 => n33, A2 => n39, ZN => ab_6_6_port);
   U57 : NOR2_X1 port map( A1 => n34, A2 => n39, ZN => ab_6_5_port);
   U58 : NOR2_X1 port map( A1 => n35, A2 => n39, ZN => ab_6_4_port);
   U59 : NOR2_X1 port map( A1 => n31, A2 => n39, ZN => ab_6_3_port);
   U60 : NOR2_X1 port map( A1 => n32, A2 => n39, ZN => ab_6_2_port);
   U61 : NOR2_X1 port map( A1 => n36, A2 => n39, ZN => ab_6_1_port);
   U62 : NOR2_X1 port map( A1 => n37, A2 => n39, ZN => ab_6_0_port);
   U63 : NOR2_X1 port map( A1 => n30, A2 => n40, ZN => ab_5_7_port);
   U64 : NOR2_X1 port map( A1 => n33, A2 => n40, ZN => ab_5_6_port);
   U65 : NOR2_X1 port map( A1 => n34, A2 => n40, ZN => ab_5_5_port);
   U66 : NOR2_X1 port map( A1 => n35, A2 => n40, ZN => ab_5_4_port);
   U67 : NOR2_X1 port map( A1 => n31, A2 => n40, ZN => ab_5_3_port);
   U68 : NOR2_X1 port map( A1 => n32, A2 => n40, ZN => ab_5_2_port);
   U69 : NOR2_X1 port map( A1 => n36, A2 => n40, ZN => ab_5_1_port);
   U70 : NOR2_X1 port map( A1 => n37, A2 => n40, ZN => ab_5_0_port);
   U71 : NOR2_X1 port map( A1 => n30, A2 => n41, ZN => ab_4_7_port);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n41, ZN => ab_4_6_port);
   U73 : NOR2_X1 port map( A1 => n34, A2 => n41, ZN => ab_4_5_port);
   U74 : NOR2_X1 port map( A1 => n35, A2 => n41, ZN => ab_4_4_port);
   U75 : NOR2_X1 port map( A1 => n31, A2 => n41, ZN => ab_4_3_port);
   U76 : NOR2_X1 port map( A1 => n32, A2 => n41, ZN => ab_4_2_port);
   U77 : NOR2_X1 port map( A1 => n36, A2 => n41, ZN => ab_4_1_port);
   U78 : NOR2_X1 port map( A1 => n37, A2 => n41, ZN => ab_4_0_port);
   U79 : NOR2_X1 port map( A1 => n30, A2 => n42, ZN => ab_3_7_port);
   U80 : NOR2_X1 port map( A1 => n33, A2 => n42, ZN => ab_3_6_port);
   U81 : NOR2_X1 port map( A1 => n34, A2 => n42, ZN => ab_3_5_port);
   U82 : NOR2_X1 port map( A1 => n35, A2 => n42, ZN => ab_3_4_port);
   U83 : NOR2_X1 port map( A1 => n31, A2 => n42, ZN => ab_3_3_port);
   U84 : NOR2_X1 port map( A1 => n32, A2 => n42, ZN => ab_3_2_port);
   U85 : NOR2_X1 port map( A1 => n36, A2 => n42, ZN => ab_3_1_port);
   U86 : NOR2_X1 port map( A1 => n37, A2 => n42, ZN => ab_3_0_port);
   U87 : NOR2_X1 port map( A1 => n30, A2 => n43, ZN => ab_2_7_port);
   U88 : NOR2_X1 port map( A1 => n33, A2 => n43, ZN => ab_2_6_port);
   U89 : NOR2_X1 port map( A1 => n34, A2 => n43, ZN => ab_2_5_port);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n43, ZN => ab_2_4_port);
   U91 : NOR2_X1 port map( A1 => n31, A2 => n43, ZN => ab_2_3_port);
   U92 : NOR2_X1 port map( A1 => n32, A2 => n43, ZN => ab_2_2_port);
   U93 : NOR2_X1 port map( A1 => n36, A2 => n43, ZN => ab_2_1_port);
   U94 : NOR2_X1 port map( A1 => n37, A2 => n43, ZN => ab_2_0_port);
   U95 : NOR2_X1 port map( A1 => n30, A2 => n44, ZN => ab_1_7_port);
   U96 : NOR2_X1 port map( A1 => n33, A2 => n44, ZN => ab_1_6_port);
   U97 : NOR2_X1 port map( A1 => n34, A2 => n44, ZN => ab_1_5_port);
   U98 : NOR2_X1 port map( A1 => n35, A2 => n44, ZN => ab_1_4_port);
   U99 : NOR2_X1 port map( A1 => n31, A2 => n44, ZN => ab_1_3_port);
   U100 : NOR2_X1 port map( A1 => n32, A2 => n44, ZN => ab_1_2_port);
   U101 : NOR2_X1 port map( A1 => n36, A2 => n44, ZN => ab_1_1_port);
   U102 : NOR2_X1 port map( A1 => n37, A2 => n44, ZN => ab_1_0_port);
   U103 : NOR2_X1 port map( A1 => n30, A2 => n45, ZN => ab_0_7_port);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n45, ZN => ab_0_6_port);
   U105 : NOR2_X1 port map( A1 => n34, A2 => n45, ZN => ab_0_5_port);
   U106 : NOR2_X1 port map( A1 => n35, A2 => n45, ZN => ab_0_4_port);
   U107 : NOR2_X1 port map( A1 => n31, A2 => n45, ZN => ab_0_3_port);
   U108 : NOR2_X1 port map( A1 => n32, A2 => n45, ZN => ab_0_2_port);
   U109 : NOR2_X1 port map( A1 => n36, A2 => n45, ZN => ab_0_1_port);
   U110 : NOR2_X1 port map( A1 => n37, A2 => n45, ZN => PRODUCT(0));
   n47 <= '0';

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_6_DW01_add_0_DW01_add_5 is

   port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (13 downto 0);  CO : out std_logic);

end shift_pow2_N8_6_DW01_add_0_DW01_add_5;

architecture SYN_cla of shift_pow2_N8_6_DW01_add_0_DW01_add_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, n1, SUM_7_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SUM <= ( SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, SUM_7_port, A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n1);
   U3 : INV_X1 port map( A => n12, ZN => n7);
   U4 : INV_X1 port map( A => n24, ZN => n4);
   U5 : INV_X1 port map( A => n27, ZN => n5);
   U6 : INV_X1 port map( A => n16, ZN => n8);
   U7 : INV_X1 port map( A => n32, ZN => n6);
   U8 : INV_X1 port map( A => n20, ZN => n3);
   U9 : XNOR2_X1 port map( A => B(13), B => n17, ZN => SUM_13_port);
   U10 : AND2_X1 port map( A1 => n16, A2 => n1, ZN => SUM_7_port);
   U11 : XNOR2_X1 port map( A => n9, B => n10, ZN => SUM_9_port);
   U12 : NOR2_X1 port map( A1 => n7, A2 => n11, ZN => n10);
   U13 : XOR2_X1 port map( A => n8, B => n13, Z => SUM_8_port);
   U14 : AND2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U15 : AOI21_X1 port map( B1 => n18, B2 => n3, A => n19, ZN => n17);
   U16 : XOR2_X1 port map( A => n18, B => n21, Z => SUM_12_port);
   U17 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U18 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n19);
   U19 : NOR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n20);
   U20 : OAI211_X1 port map( C1 => n22, C2 => n23, A => n24, B => n25, ZN => 
                           n18);
   U21 : OR4_X1 port map( A1 => n26, A2 => n27, A3 => n23, A4 => n11, ZN => n25
                           );
   U22 : AOI21_X1 port map( B1 => n5, B2 => n28, A => n6, ZN => n22);
   U23 : OAI21_X1 port map( B1 => n11, B2 => n15, A => n12, ZN => n28);
   U24 : XNOR2_X1 port map( A => n29, B => n30, ZN => SUM_11_port);
   U25 : NOR2_X1 port map( A1 => n23, A2 => n4, ZN => n30);
   U26 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n24);
   U27 : NOR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n23);
   U28 : AOI21_X1 port map( B1 => n31, B2 => n5, A => n6, ZN => n29);
   U29 : XNOR2_X1 port map( A => n33, B => n31, ZN => SUM_10_port);
   U30 : OAI21_X1 port map( B1 => n11, B2 => n9, A => n12, ZN => n31);
   U31 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n12);
   U32 : AND2_X1 port map( A1 => n26, A2 => n15, ZN => n9);
   U33 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n15);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n14, ZN => n26);
   U35 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n14);
   U36 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n16);
   U37 : NOR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n11);
   U38 : NAND2_X1 port map( A1 => n32, A2 => n5, ZN => n33);
   U39 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n27);
   U40 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n32);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_6_DW02_mult_0_DW02_mult_5 is

   port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  PRODUCT 
         : out std_logic_vector (15 downto 0));

end shift_pow2_N8_6_DW02_mult_0_DW02_mult_5;

architecture SYN_csa of shift_pow2_N8_6_DW02_mult_0_DW02_mult_5 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component shift_pow2_N8_6_DW01_add_0_DW01_add_5
      port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (13 downto 0);  CO : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, ab_7_4_port, 
      ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_7_port, ab_3_6_port, 
      ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, 
      ab_3_0_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, ab_2_4_port, 
      ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, ab_1_7_port, 
      ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_2_port, 
      ab_1_1_port, ab_1_0_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, 
      SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, SUMB_7_0_port, SUMB_6_6_port
      , SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, 
      SUMB_6_1_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_6_port, SUMB_4_5_port, 
      SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_6_port
      , SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, 
      SUMB_3_1_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n_1035 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => 
                           SUMB_7_0_port);
   S4_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S4_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S4_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S4_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S4_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S5_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           ab_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S3_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           ab_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S3_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           ab_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S3_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           ab_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S3_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           ab_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n7, CI => n13, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n6, CI => n14, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n5, CI => n12, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n4, CI => n11, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n3, CI => n10, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n2, CI => n9, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S3_2_6 : FA_X1 port map( A => ab_2_6_port, B => n8, CI => ab_1_7_port, CO =>
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   FS_1 : shift_pow2_N8_6_DW01_add_0_DW01_add_5 port map( A(13) => n46, A(12) 
                           => n18, A(11) => n21, A(10) => n19, A(9) => n22, 
                           A(8) => n27, A(7) => n20, A(6) => n17, A(5) => 
                           SUMB_7_0_port, A(4) => A1_4_port, A(3) => A1_3_port,
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(13) => n15, B(12) => n29, B(11) => n26,
                           B(10) => n25, B(9) => n24, B(8) => n28, B(7) => n23,
                           B(6) => n46, B(5) => n47, B(4) => n47, B(3) => n47, 
                           B(2) => n47, B(1) => n47, B(0) => X_Logic0_port, CI 
                           => X_Logic0_port, SUM(13) => PRODUCT(15), SUM(12) =>
                           PRODUCT(14), SUM(11) => PRODUCT(13), SUM(10) => 
                           PRODUCT(12), SUM(9) => PRODUCT(11), SUM(8) => 
                           PRODUCT(10), SUM(7) => PRODUCT(9), SUM(6) => 
                           PRODUCT(8), SUM(5) => PRODUCT(7), SUM(4) => 
                           PRODUCT(6), SUM(3) => PRODUCT(5), SUM(2) => 
                           PRODUCT(4), SUM(1) => PRODUCT(3), SUM(0) => 
                           PRODUCT(2), CO => n_1035);
   U2 : INV_X1 port map( A => B(4), ZN => n35);
   U3 : INV_X1 port map( A => B(5), ZN => n34);
   U4 : INV_X1 port map( A => B(6), ZN => n33);
   U5 : INV_X1 port map( A => B(7), ZN => n30);
   U6 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n2);
   U7 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n3);
   U8 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n4);
   U9 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n5);
   U10 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n6);
   U11 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n7);
   U12 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n8);
   U13 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n9);
   U14 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n10);
   U15 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n11);
   U16 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n12);
   U17 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n13);
   U18 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n14);
   U19 : AND2_X1 port map( A1 => CARRYB_7_6_port, A2 => ab_7_7_port, ZN => n15)
                           ;
   U20 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U21 : XOR2_X1 port map( A => CARRYB_7_0_port, B => SUMB_7_1_port, Z => n17);
   U22 : XOR2_X1 port map( A => CARRYB_7_6_port, B => ab_7_7_port, Z => n18);
   U23 : XOR2_X1 port map( A => CARRYB_7_4_port, B => SUMB_7_5_port, Z => n19);
   U24 : XOR2_X1 port map( A => CARRYB_7_1_port, B => SUMB_7_2_port, Z => n20);
   U25 : XOR2_X1 port map( A => CARRYB_7_5_port, B => SUMB_7_6_port, Z => n21);
   U26 : XOR2_X1 port map( A => CARRYB_7_3_port, B => SUMB_7_4_port, Z => n22);
   U27 : AND2_X1 port map( A1 => CARRYB_7_0_port, A2 => SUMB_7_1_port, ZN => 
                           n23);
   U28 : AND2_X1 port map( A1 => CARRYB_7_2_port, A2 => SUMB_7_3_port, ZN => 
                           n24);
   U29 : AND2_X1 port map( A1 => CARRYB_7_3_port, A2 => SUMB_7_4_port, ZN => 
                           n25);
   U30 : AND2_X1 port map( A1 => CARRYB_7_4_port, A2 => SUMB_7_5_port, ZN => 
                           n26);
   U31 : XOR2_X1 port map( A => CARRYB_7_2_port, B => SUMB_7_3_port, Z => n27);
   U32 : AND2_X1 port map( A1 => CARRYB_7_1_port, A2 => SUMB_7_2_port, ZN => 
                           n28);
   U33 : AND2_X1 port map( A1 => CARRYB_7_5_port, A2 => SUMB_7_6_port, ZN => 
                           n29);
   U34 : INV_X1 port map( A => B(3), ZN => n31);
   U35 : INV_X1 port map( A => B(2), ZN => n32);
   U36 : INV_X1 port map( A => B(1), ZN => n36);
   U37 : INV_X1 port map( A => B(0), ZN => n37);
   U38 : INV_X1 port map( A => A(7), ZN => n38);
   U39 : INV_X1 port map( A => A(0), ZN => n45);
   U40 : INV_X1 port map( A => A(1), ZN => n44);
   U41 : INV_X1 port map( A => A(3), ZN => n42);
   U42 : INV_X1 port map( A => A(4), ZN => n41);
   U43 : INV_X1 port map( A => A(5), ZN => n40);
   U44 : INV_X1 port map( A => A(6), ZN => n39);
   U45 : INV_X1 port map( A => A(2), ZN => n43);
   n46 <= '0';
   U47 : NOR2_X1 port map( A1 => n38, A2 => n30, ZN => ab_7_7_port);
   U48 : NOR2_X1 port map( A1 => n38, A2 => n33, ZN => ab_7_6_port);
   U49 : NOR2_X1 port map( A1 => n38, A2 => n34, ZN => ab_7_5_port);
   U50 : NOR2_X1 port map( A1 => n38, A2 => n35, ZN => ab_7_4_port);
   U51 : NOR2_X1 port map( A1 => n38, A2 => n31, ZN => ab_7_3_port);
   U52 : NOR2_X1 port map( A1 => n38, A2 => n32, ZN => ab_7_2_port);
   U53 : NOR2_X1 port map( A1 => n38, A2 => n36, ZN => ab_7_1_port);
   U54 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => ab_7_0_port);
   U55 : NOR2_X1 port map( A1 => n30, A2 => n39, ZN => ab_6_7_port);
   U56 : NOR2_X1 port map( A1 => n33, A2 => n39, ZN => ab_6_6_port);
   U57 : NOR2_X1 port map( A1 => n34, A2 => n39, ZN => ab_6_5_port);
   U58 : NOR2_X1 port map( A1 => n35, A2 => n39, ZN => ab_6_4_port);
   U59 : NOR2_X1 port map( A1 => n31, A2 => n39, ZN => ab_6_3_port);
   U60 : NOR2_X1 port map( A1 => n32, A2 => n39, ZN => ab_6_2_port);
   U61 : NOR2_X1 port map( A1 => n36, A2 => n39, ZN => ab_6_1_port);
   U62 : NOR2_X1 port map( A1 => n37, A2 => n39, ZN => ab_6_0_port);
   U63 : NOR2_X1 port map( A1 => n30, A2 => n40, ZN => ab_5_7_port);
   U64 : NOR2_X1 port map( A1 => n33, A2 => n40, ZN => ab_5_6_port);
   U65 : NOR2_X1 port map( A1 => n34, A2 => n40, ZN => ab_5_5_port);
   U66 : NOR2_X1 port map( A1 => n35, A2 => n40, ZN => ab_5_4_port);
   U67 : NOR2_X1 port map( A1 => n31, A2 => n40, ZN => ab_5_3_port);
   U68 : NOR2_X1 port map( A1 => n32, A2 => n40, ZN => ab_5_2_port);
   U69 : NOR2_X1 port map( A1 => n36, A2 => n40, ZN => ab_5_1_port);
   U70 : NOR2_X1 port map( A1 => n37, A2 => n40, ZN => ab_5_0_port);
   U71 : NOR2_X1 port map( A1 => n30, A2 => n41, ZN => ab_4_7_port);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n41, ZN => ab_4_6_port);
   U73 : NOR2_X1 port map( A1 => n34, A2 => n41, ZN => ab_4_5_port);
   U74 : NOR2_X1 port map( A1 => n35, A2 => n41, ZN => ab_4_4_port);
   U75 : NOR2_X1 port map( A1 => n31, A2 => n41, ZN => ab_4_3_port);
   U76 : NOR2_X1 port map( A1 => n32, A2 => n41, ZN => ab_4_2_port);
   U77 : NOR2_X1 port map( A1 => n36, A2 => n41, ZN => ab_4_1_port);
   U78 : NOR2_X1 port map( A1 => n37, A2 => n41, ZN => ab_4_0_port);
   U79 : NOR2_X1 port map( A1 => n30, A2 => n42, ZN => ab_3_7_port);
   U80 : NOR2_X1 port map( A1 => n33, A2 => n42, ZN => ab_3_6_port);
   U81 : NOR2_X1 port map( A1 => n34, A2 => n42, ZN => ab_3_5_port);
   U82 : NOR2_X1 port map( A1 => n35, A2 => n42, ZN => ab_3_4_port);
   U83 : NOR2_X1 port map( A1 => n31, A2 => n42, ZN => ab_3_3_port);
   U84 : NOR2_X1 port map( A1 => n32, A2 => n42, ZN => ab_3_2_port);
   U85 : NOR2_X1 port map( A1 => n36, A2 => n42, ZN => ab_3_1_port);
   U86 : NOR2_X1 port map( A1 => n37, A2 => n42, ZN => ab_3_0_port);
   U87 : NOR2_X1 port map( A1 => n30, A2 => n43, ZN => ab_2_7_port);
   U88 : NOR2_X1 port map( A1 => n33, A2 => n43, ZN => ab_2_6_port);
   U89 : NOR2_X1 port map( A1 => n34, A2 => n43, ZN => ab_2_5_port);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n43, ZN => ab_2_4_port);
   U91 : NOR2_X1 port map( A1 => n31, A2 => n43, ZN => ab_2_3_port);
   U92 : NOR2_X1 port map( A1 => n32, A2 => n43, ZN => ab_2_2_port);
   U93 : NOR2_X1 port map( A1 => n36, A2 => n43, ZN => ab_2_1_port);
   U94 : NOR2_X1 port map( A1 => n37, A2 => n43, ZN => ab_2_0_port);
   U95 : NOR2_X1 port map( A1 => n30, A2 => n44, ZN => ab_1_7_port);
   U96 : NOR2_X1 port map( A1 => n33, A2 => n44, ZN => ab_1_6_port);
   U97 : NOR2_X1 port map( A1 => n34, A2 => n44, ZN => ab_1_5_port);
   U98 : NOR2_X1 port map( A1 => n35, A2 => n44, ZN => ab_1_4_port);
   U99 : NOR2_X1 port map( A1 => n31, A2 => n44, ZN => ab_1_3_port);
   U100 : NOR2_X1 port map( A1 => n32, A2 => n44, ZN => ab_1_2_port);
   U101 : NOR2_X1 port map( A1 => n36, A2 => n44, ZN => ab_1_1_port);
   U102 : NOR2_X1 port map( A1 => n37, A2 => n44, ZN => ab_1_0_port);
   U103 : NOR2_X1 port map( A1 => n30, A2 => n45, ZN => ab_0_7_port);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n45, ZN => ab_0_6_port);
   U105 : NOR2_X1 port map( A1 => n34, A2 => n45, ZN => ab_0_5_port);
   U106 : NOR2_X1 port map( A1 => n35, A2 => n45, ZN => ab_0_4_port);
   U107 : NOR2_X1 port map( A1 => n31, A2 => n45, ZN => ab_0_3_port);
   U108 : NOR2_X1 port map( A1 => n32, A2 => n45, ZN => ab_0_2_port);
   U109 : NOR2_X1 port map( A1 => n36, A2 => n45, ZN => ab_0_1_port);
   U110 : NOR2_X1 port map( A1 => n37, A2 => n45, ZN => PRODUCT(0));
   n47 <= '0';

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_5_DW01_add_0_DW01_add_4 is

   port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (13 downto 0);  CO : out std_logic);

end shift_pow2_N8_5_DW01_add_0_DW01_add_4;

architecture SYN_cla of shift_pow2_N8_5_DW01_add_0_DW01_add_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, n1, SUM_7_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SUM <= ( SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, SUM_7_port, A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n1);
   U3 : INV_X1 port map( A => n12, ZN => n7);
   U4 : INV_X1 port map( A => n24, ZN => n4);
   U5 : INV_X1 port map( A => n27, ZN => n5);
   U6 : INV_X1 port map( A => n16, ZN => n8);
   U7 : INV_X1 port map( A => n32, ZN => n6);
   U8 : INV_X1 port map( A => n20, ZN => n3);
   U9 : XNOR2_X1 port map( A => B(13), B => n17, ZN => SUM_13_port);
   U10 : AND2_X1 port map( A1 => n16, A2 => n1, ZN => SUM_7_port);
   U11 : XNOR2_X1 port map( A => n9, B => n10, ZN => SUM_9_port);
   U12 : NOR2_X1 port map( A1 => n7, A2 => n11, ZN => n10);
   U13 : XOR2_X1 port map( A => n8, B => n13, Z => SUM_8_port);
   U14 : AND2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U15 : AOI21_X1 port map( B1 => n18, B2 => n3, A => n19, ZN => n17);
   U16 : XOR2_X1 port map( A => n18, B => n21, Z => SUM_12_port);
   U17 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U18 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n19);
   U19 : NOR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n20);
   U20 : OAI211_X1 port map( C1 => n22, C2 => n23, A => n24, B => n25, ZN => 
                           n18);
   U21 : OR4_X1 port map( A1 => n26, A2 => n27, A3 => n23, A4 => n11, ZN => n25
                           );
   U22 : AOI21_X1 port map( B1 => n5, B2 => n28, A => n6, ZN => n22);
   U23 : OAI21_X1 port map( B1 => n11, B2 => n15, A => n12, ZN => n28);
   U24 : XNOR2_X1 port map( A => n29, B => n30, ZN => SUM_11_port);
   U25 : NOR2_X1 port map( A1 => n23, A2 => n4, ZN => n30);
   U26 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n24);
   U27 : NOR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n23);
   U28 : AOI21_X1 port map( B1 => n31, B2 => n5, A => n6, ZN => n29);
   U29 : XNOR2_X1 port map( A => n33, B => n31, ZN => SUM_10_port);
   U30 : OAI21_X1 port map( B1 => n11, B2 => n9, A => n12, ZN => n31);
   U31 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n12);
   U32 : AND2_X1 port map( A1 => n26, A2 => n15, ZN => n9);
   U33 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n15);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n14, ZN => n26);
   U35 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n14);
   U36 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n16);
   U37 : NOR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n11);
   U38 : NAND2_X1 port map( A1 => n32, A2 => n5, ZN => n33);
   U39 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n27);
   U40 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n32);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_5_DW02_mult_0_DW02_mult_4 is

   port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  PRODUCT 
         : out std_logic_vector (15 downto 0));

end shift_pow2_N8_5_DW02_mult_0_DW02_mult_4;

architecture SYN_csa of shift_pow2_N8_5_DW02_mult_0_DW02_mult_4 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component shift_pow2_N8_5_DW01_add_0_DW01_add_4
      port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (13 downto 0);  CO : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, ab_7_4_port, 
      ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_7_port, ab_3_6_port, 
      ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, 
      ab_3_0_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, ab_2_4_port, 
      ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, ab_1_7_port, 
      ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_2_port, 
      ab_1_1_port, ab_1_0_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, 
      SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, SUMB_7_0_port, SUMB_6_6_port
      , SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, 
      SUMB_6_1_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_6_port, SUMB_4_5_port, 
      SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_6_port
      , SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, 
      SUMB_3_1_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n_1047 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => 
                           SUMB_7_0_port);
   S4_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S4_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S4_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S4_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S4_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S5_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           ab_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S3_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           ab_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S3_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           ab_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S3_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           ab_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S3_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           ab_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n7, CI => n13, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n6, CI => n12, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n5, CI => n14, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n4, CI => n11, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n3, CI => n10, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n2, CI => n9, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S3_2_6 : FA_X1 port map( A => ab_2_6_port, B => n8, CI => ab_1_7_port, CO =>
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   FS_1 : shift_pow2_N8_5_DW01_add_0_DW01_add_4 port map( A(13) => n46, A(12) 
                           => n17, A(11) => n20, A(10) => n19, A(9) => n21, 
                           A(8) => n27, A(7) => n22, A(6) => n18, A(5) => 
                           SUMB_7_0_port, A(4) => A1_4_port, A(3) => A1_3_port,
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(13) => n15, B(12) => n29, B(11) => n26,
                           B(10) => n23, B(9) => n25, B(8) => n28, B(7) => n24,
                           B(6) => n46, B(5) => n47, B(4) => n47, B(3) => n47, 
                           B(2) => n47, B(1) => n47, B(0) => X_Logic0_port, CI 
                           => X_Logic0_port, SUM(13) => PRODUCT(15), SUM(12) =>
                           PRODUCT(14), SUM(11) => PRODUCT(13), SUM(10) => 
                           PRODUCT(12), SUM(9) => PRODUCT(11), SUM(8) => 
                           PRODUCT(10), SUM(7) => PRODUCT(9), SUM(6) => 
                           PRODUCT(8), SUM(5) => PRODUCT(7), SUM(4) => 
                           PRODUCT(6), SUM(3) => PRODUCT(5), SUM(2) => 
                           PRODUCT(4), SUM(1) => PRODUCT(3), SUM(0) => 
                           PRODUCT(2), CO => n_1047);
   U2 : INV_X1 port map( A => B(4), ZN => n35);
   U3 : INV_X1 port map( A => B(5), ZN => n34);
   U4 : INV_X1 port map( A => B(6), ZN => n33);
   U5 : INV_X1 port map( A => B(7), ZN => n30);
   U6 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n2);
   U7 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n3);
   U8 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n4);
   U9 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n5);
   U10 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n6);
   U11 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n7);
   U12 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n8);
   U13 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n9);
   U14 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n10);
   U15 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n11);
   U16 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n12);
   U17 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n13);
   U18 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n14);
   U19 : AND2_X1 port map( A1 => CARRYB_7_6_port, A2 => ab_7_7_port, ZN => n15)
                           ;
   U20 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U21 : XOR2_X1 port map( A => CARRYB_7_6_port, B => ab_7_7_port, Z => n17);
   U22 : XOR2_X1 port map( A => CARRYB_7_0_port, B => SUMB_7_1_port, Z => n18);
   U23 : XOR2_X1 port map( A => CARRYB_7_4_port, B => SUMB_7_5_port, Z => n19);
   U24 : XOR2_X1 port map( A => CARRYB_7_5_port, B => SUMB_7_6_port, Z => n20);
   U25 : XOR2_X1 port map( A => CARRYB_7_3_port, B => SUMB_7_4_port, Z => n21);
   U26 : XOR2_X1 port map( A => CARRYB_7_1_port, B => SUMB_7_2_port, Z => n22);
   U27 : AND2_X1 port map( A1 => CARRYB_7_3_port, A2 => SUMB_7_4_port, ZN => 
                           n23);
   U28 : AND2_X1 port map( A1 => CARRYB_7_0_port, A2 => SUMB_7_1_port, ZN => 
                           n24);
   U29 : AND2_X1 port map( A1 => CARRYB_7_2_port, A2 => SUMB_7_3_port, ZN => 
                           n25);
   U30 : AND2_X1 port map( A1 => CARRYB_7_4_port, A2 => SUMB_7_5_port, ZN => 
                           n26);
   U31 : XOR2_X1 port map( A => CARRYB_7_2_port, B => SUMB_7_3_port, Z => n27);
   U32 : AND2_X1 port map( A1 => CARRYB_7_1_port, A2 => SUMB_7_2_port, ZN => 
                           n28);
   U33 : AND2_X1 port map( A1 => CARRYB_7_5_port, A2 => SUMB_7_6_port, ZN => 
                           n29);
   U34 : INV_X1 port map( A => B(3), ZN => n31);
   U35 : INV_X1 port map( A => B(2), ZN => n32);
   U36 : INV_X1 port map( A => B(1), ZN => n36);
   U37 : INV_X1 port map( A => B(0), ZN => n37);
   U38 : INV_X1 port map( A => A(7), ZN => n38);
   U39 : INV_X1 port map( A => A(0), ZN => n45);
   U40 : INV_X1 port map( A => A(1), ZN => n44);
   U41 : INV_X1 port map( A => A(3), ZN => n42);
   U42 : INV_X1 port map( A => A(2), ZN => n43);
   U43 : INV_X1 port map( A => A(4), ZN => n41);
   U44 : INV_X1 port map( A => A(5), ZN => n40);
   U45 : INV_X1 port map( A => A(6), ZN => n39);
   n46 <= '0';
   U47 : NOR2_X1 port map( A1 => n38, A2 => n30, ZN => ab_7_7_port);
   U48 : NOR2_X1 port map( A1 => n38, A2 => n33, ZN => ab_7_6_port);
   U49 : NOR2_X1 port map( A1 => n38, A2 => n34, ZN => ab_7_5_port);
   U50 : NOR2_X1 port map( A1 => n38, A2 => n35, ZN => ab_7_4_port);
   U51 : NOR2_X1 port map( A1 => n38, A2 => n31, ZN => ab_7_3_port);
   U52 : NOR2_X1 port map( A1 => n38, A2 => n32, ZN => ab_7_2_port);
   U53 : NOR2_X1 port map( A1 => n38, A2 => n36, ZN => ab_7_1_port);
   U54 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => ab_7_0_port);
   U55 : NOR2_X1 port map( A1 => n30, A2 => n39, ZN => ab_6_7_port);
   U56 : NOR2_X1 port map( A1 => n33, A2 => n39, ZN => ab_6_6_port);
   U57 : NOR2_X1 port map( A1 => n34, A2 => n39, ZN => ab_6_5_port);
   U58 : NOR2_X1 port map( A1 => n35, A2 => n39, ZN => ab_6_4_port);
   U59 : NOR2_X1 port map( A1 => n31, A2 => n39, ZN => ab_6_3_port);
   U60 : NOR2_X1 port map( A1 => n32, A2 => n39, ZN => ab_6_2_port);
   U61 : NOR2_X1 port map( A1 => n36, A2 => n39, ZN => ab_6_1_port);
   U62 : NOR2_X1 port map( A1 => n37, A2 => n39, ZN => ab_6_0_port);
   U63 : NOR2_X1 port map( A1 => n30, A2 => n40, ZN => ab_5_7_port);
   U64 : NOR2_X1 port map( A1 => n33, A2 => n40, ZN => ab_5_6_port);
   U65 : NOR2_X1 port map( A1 => n34, A2 => n40, ZN => ab_5_5_port);
   U66 : NOR2_X1 port map( A1 => n35, A2 => n40, ZN => ab_5_4_port);
   U67 : NOR2_X1 port map( A1 => n31, A2 => n40, ZN => ab_5_3_port);
   U68 : NOR2_X1 port map( A1 => n32, A2 => n40, ZN => ab_5_2_port);
   U69 : NOR2_X1 port map( A1 => n36, A2 => n40, ZN => ab_5_1_port);
   U70 : NOR2_X1 port map( A1 => n37, A2 => n40, ZN => ab_5_0_port);
   U71 : NOR2_X1 port map( A1 => n30, A2 => n41, ZN => ab_4_7_port);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n41, ZN => ab_4_6_port);
   U73 : NOR2_X1 port map( A1 => n34, A2 => n41, ZN => ab_4_5_port);
   U74 : NOR2_X1 port map( A1 => n35, A2 => n41, ZN => ab_4_4_port);
   U75 : NOR2_X1 port map( A1 => n31, A2 => n41, ZN => ab_4_3_port);
   U76 : NOR2_X1 port map( A1 => n32, A2 => n41, ZN => ab_4_2_port);
   U77 : NOR2_X1 port map( A1 => n36, A2 => n41, ZN => ab_4_1_port);
   U78 : NOR2_X1 port map( A1 => n37, A2 => n41, ZN => ab_4_0_port);
   U79 : NOR2_X1 port map( A1 => n30, A2 => n42, ZN => ab_3_7_port);
   U80 : NOR2_X1 port map( A1 => n33, A2 => n42, ZN => ab_3_6_port);
   U81 : NOR2_X1 port map( A1 => n34, A2 => n42, ZN => ab_3_5_port);
   U82 : NOR2_X1 port map( A1 => n35, A2 => n42, ZN => ab_3_4_port);
   U83 : NOR2_X1 port map( A1 => n31, A2 => n42, ZN => ab_3_3_port);
   U84 : NOR2_X1 port map( A1 => n32, A2 => n42, ZN => ab_3_2_port);
   U85 : NOR2_X1 port map( A1 => n36, A2 => n42, ZN => ab_3_1_port);
   U86 : NOR2_X1 port map( A1 => n37, A2 => n42, ZN => ab_3_0_port);
   U87 : NOR2_X1 port map( A1 => n30, A2 => n43, ZN => ab_2_7_port);
   U88 : NOR2_X1 port map( A1 => n33, A2 => n43, ZN => ab_2_6_port);
   U89 : NOR2_X1 port map( A1 => n34, A2 => n43, ZN => ab_2_5_port);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n43, ZN => ab_2_4_port);
   U91 : NOR2_X1 port map( A1 => n31, A2 => n43, ZN => ab_2_3_port);
   U92 : NOR2_X1 port map( A1 => n32, A2 => n43, ZN => ab_2_2_port);
   U93 : NOR2_X1 port map( A1 => n36, A2 => n43, ZN => ab_2_1_port);
   U94 : NOR2_X1 port map( A1 => n37, A2 => n43, ZN => ab_2_0_port);
   U95 : NOR2_X1 port map( A1 => n30, A2 => n44, ZN => ab_1_7_port);
   U96 : NOR2_X1 port map( A1 => n33, A2 => n44, ZN => ab_1_6_port);
   U97 : NOR2_X1 port map( A1 => n34, A2 => n44, ZN => ab_1_5_port);
   U98 : NOR2_X1 port map( A1 => n35, A2 => n44, ZN => ab_1_4_port);
   U99 : NOR2_X1 port map( A1 => n31, A2 => n44, ZN => ab_1_3_port);
   U100 : NOR2_X1 port map( A1 => n32, A2 => n44, ZN => ab_1_2_port);
   U101 : NOR2_X1 port map( A1 => n36, A2 => n44, ZN => ab_1_1_port);
   U102 : NOR2_X1 port map( A1 => n37, A2 => n44, ZN => ab_1_0_port);
   U103 : NOR2_X1 port map( A1 => n30, A2 => n45, ZN => ab_0_7_port);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n45, ZN => ab_0_6_port);
   U105 : NOR2_X1 port map( A1 => n34, A2 => n45, ZN => ab_0_5_port);
   U106 : NOR2_X1 port map( A1 => n35, A2 => n45, ZN => ab_0_4_port);
   U107 : NOR2_X1 port map( A1 => n31, A2 => n45, ZN => ab_0_3_port);
   U108 : NOR2_X1 port map( A1 => n32, A2 => n45, ZN => ab_0_2_port);
   U109 : NOR2_X1 port map( A1 => n36, A2 => n45, ZN => ab_0_1_port);
   U110 : NOR2_X1 port map( A1 => n37, A2 => n45, ZN => PRODUCT(0));
   n47 <= '0';

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_4_DW01_add_0_DW01_add_3 is

   port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (13 downto 0);  CO : out std_logic);

end shift_pow2_N8_4_DW01_add_0_DW01_add_3;

architecture SYN_cla of shift_pow2_N8_4_DW01_add_0_DW01_add_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, n1, SUM_7_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SUM <= ( SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, SUM_7_port, A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n1);
   U3 : INV_X1 port map( A => n24, ZN => n4);
   U4 : INV_X1 port map( A => n12, ZN => n7);
   U5 : INV_X1 port map( A => n27, ZN => n5);
   U6 : INV_X1 port map( A => n16, ZN => n8);
   U7 : INV_X1 port map( A => n32, ZN => n6);
   U8 : INV_X1 port map( A => n20, ZN => n3);
   U9 : XNOR2_X1 port map( A => B(13), B => n17, ZN => SUM_13_port);
   U10 : AND2_X1 port map( A1 => n16, A2 => n1, ZN => SUM_7_port);
   U11 : XNOR2_X1 port map( A => n9, B => n10, ZN => SUM_9_port);
   U12 : NOR2_X1 port map( A1 => n7, A2 => n11, ZN => n10);
   U13 : XOR2_X1 port map( A => n8, B => n13, Z => SUM_8_port);
   U14 : AND2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U15 : AOI21_X1 port map( B1 => n18, B2 => n3, A => n19, ZN => n17);
   U16 : XOR2_X1 port map( A => n18, B => n21, Z => SUM_12_port);
   U17 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U18 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n19);
   U19 : NOR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n20);
   U20 : OAI211_X1 port map( C1 => n22, C2 => n23, A => n24, B => n25, ZN => 
                           n18);
   U21 : OR4_X1 port map( A1 => n26, A2 => n27, A3 => n23, A4 => n11, ZN => n25
                           );
   U22 : AOI21_X1 port map( B1 => n5, B2 => n28, A => n6, ZN => n22);
   U23 : OAI21_X1 port map( B1 => n11, B2 => n15, A => n12, ZN => n28);
   U24 : XNOR2_X1 port map( A => n29, B => n30, ZN => SUM_11_port);
   U25 : NOR2_X1 port map( A1 => n23, A2 => n4, ZN => n30);
   U26 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n24);
   U27 : NOR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n23);
   U28 : AOI21_X1 port map( B1 => n31, B2 => n5, A => n6, ZN => n29);
   U29 : XNOR2_X1 port map( A => n33, B => n31, ZN => SUM_10_port);
   U30 : OAI21_X1 port map( B1 => n11, B2 => n9, A => n12, ZN => n31);
   U31 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n12);
   U32 : AND2_X1 port map( A1 => n26, A2 => n15, ZN => n9);
   U33 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n15);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n14, ZN => n26);
   U35 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n14);
   U36 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n16);
   U37 : NOR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n11);
   U38 : NAND2_X1 port map( A1 => n32, A2 => n5, ZN => n33);
   U39 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n27);
   U40 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n32);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_4_DW02_mult_0_DW02_mult_3 is

   port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  PRODUCT 
         : out std_logic_vector (15 downto 0));

end shift_pow2_N8_4_DW02_mult_0_DW02_mult_3;

architecture SYN_csa of shift_pow2_N8_4_DW02_mult_0_DW02_mult_3 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component shift_pow2_N8_4_DW01_add_0_DW01_add_3
      port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (13 downto 0);  CO : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, ab_7_4_port, 
      ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_7_port, ab_3_6_port, 
      ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, 
      ab_3_0_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, ab_2_4_port, 
      ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, ab_1_7_port, 
      ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_2_port, 
      ab_1_1_port, ab_1_0_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, 
      SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, SUMB_7_0_port, SUMB_6_6_port
      , SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, 
      SUMB_6_1_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_6_port, SUMB_4_5_port, 
      SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_6_port
      , SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, 
      SUMB_3_1_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n_1059 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => 
                           SUMB_7_0_port);
   S4_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S4_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S4_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S4_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S4_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S5_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           ab_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S3_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           ab_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S3_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           ab_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S3_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           ab_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S3_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           ab_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n7, CI => n13, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n6, CI => n12, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n5, CI => n11, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n4, CI => n14, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n3, CI => n10, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n2, CI => n9, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S3_2_6 : FA_X1 port map( A => ab_2_6_port, B => n8, CI => ab_1_7_port, CO =>
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   FS_1 : shift_pow2_N8_4_DW01_add_0_DW01_add_3 port map( A(13) => n46, A(12) 
                           => n18, A(11) => n20, A(10) => n19, A(9) => n21, 
                           A(8) => n27, A(7) => n22, A(6) => n17, A(5) => 
                           SUMB_7_0_port, A(4) => A1_4_port, A(3) => A1_3_port,
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(13) => n15, B(12) => n29, B(11) => n25,
                           B(10) => n24, B(9) => n26, B(8) => n28, B(7) => n23,
                           B(6) => n46, B(5) => n47, B(4) => n47, B(3) => n47, 
                           B(2) => n47, B(1) => n47, B(0) => X_Logic0_port, CI 
                           => X_Logic0_port, SUM(13) => PRODUCT(15), SUM(12) =>
                           PRODUCT(14), SUM(11) => PRODUCT(13), SUM(10) => 
                           PRODUCT(12), SUM(9) => PRODUCT(11), SUM(8) => 
                           PRODUCT(10), SUM(7) => PRODUCT(9), SUM(6) => 
                           PRODUCT(8), SUM(5) => PRODUCT(7), SUM(4) => 
                           PRODUCT(6), SUM(3) => PRODUCT(5), SUM(2) => 
                           PRODUCT(4), SUM(1) => PRODUCT(3), SUM(0) => 
                           PRODUCT(2), CO => n_1059);
   U2 : INV_X1 port map( A => B(4), ZN => n35);
   U3 : INV_X1 port map( A => B(5), ZN => n34);
   U4 : INV_X1 port map( A => B(6), ZN => n33);
   U5 : INV_X1 port map( A => B(7), ZN => n30);
   U6 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n2);
   U7 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n3);
   U8 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n4);
   U9 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n5);
   U10 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n6);
   U11 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n7);
   U12 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n8);
   U13 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n9);
   U14 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n10);
   U15 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n11);
   U16 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n12);
   U17 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n13);
   U18 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n14);
   U19 : AND2_X1 port map( A1 => CARRYB_7_6_port, A2 => ab_7_7_port, ZN => n15)
                           ;
   U20 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U21 : XOR2_X1 port map( A => CARRYB_7_0_port, B => SUMB_7_1_port, Z => n17);
   U22 : XOR2_X1 port map( A => CARRYB_7_6_port, B => ab_7_7_port, Z => n18);
   U23 : XOR2_X1 port map( A => CARRYB_7_4_port, B => SUMB_7_5_port, Z => n19);
   U24 : XOR2_X1 port map( A => CARRYB_7_5_port, B => SUMB_7_6_port, Z => n20);
   U25 : XOR2_X1 port map( A => CARRYB_7_3_port, B => SUMB_7_4_port, Z => n21);
   U26 : XOR2_X1 port map( A => CARRYB_7_1_port, B => SUMB_7_2_port, Z => n22);
   U27 : AND2_X1 port map( A1 => CARRYB_7_0_port, A2 => SUMB_7_1_port, ZN => 
                           n23);
   U28 : AND2_X1 port map( A1 => CARRYB_7_3_port, A2 => SUMB_7_4_port, ZN => 
                           n24);
   U29 : AND2_X1 port map( A1 => CARRYB_7_4_port, A2 => SUMB_7_5_port, ZN => 
                           n25);
   U30 : AND2_X1 port map( A1 => CARRYB_7_2_port, A2 => SUMB_7_3_port, ZN => 
                           n26);
   U31 : XOR2_X1 port map( A => CARRYB_7_2_port, B => SUMB_7_3_port, Z => n27);
   U32 : AND2_X1 port map( A1 => CARRYB_7_1_port, A2 => SUMB_7_2_port, ZN => 
                           n28);
   U33 : AND2_X1 port map( A1 => CARRYB_7_5_port, A2 => SUMB_7_6_port, ZN => 
                           n29);
   U34 : INV_X1 port map( A => B(2), ZN => n32);
   U35 : INV_X1 port map( A => B(1), ZN => n36);
   U36 : INV_X1 port map( A => B(3), ZN => n31);
   U37 : INV_X1 port map( A => B(0), ZN => n37);
   U38 : INV_X1 port map( A => A(7), ZN => n38);
   U39 : INV_X1 port map( A => A(0), ZN => n45);
   U40 : INV_X1 port map( A => A(1), ZN => n44);
   U41 : INV_X1 port map( A => A(3), ZN => n42);
   U42 : INV_X1 port map( A => A(4), ZN => n41);
   U43 : INV_X1 port map( A => A(5), ZN => n40);
   U44 : INV_X1 port map( A => A(6), ZN => n39);
   U45 : INV_X1 port map( A => A(2), ZN => n43);
   n46 <= '0';
   U47 : NOR2_X1 port map( A1 => n38, A2 => n30, ZN => ab_7_7_port);
   U48 : NOR2_X1 port map( A1 => n38, A2 => n33, ZN => ab_7_6_port);
   U49 : NOR2_X1 port map( A1 => n38, A2 => n34, ZN => ab_7_5_port);
   U50 : NOR2_X1 port map( A1 => n38, A2 => n35, ZN => ab_7_4_port);
   U51 : NOR2_X1 port map( A1 => n38, A2 => n31, ZN => ab_7_3_port);
   U52 : NOR2_X1 port map( A1 => n38, A2 => n32, ZN => ab_7_2_port);
   U53 : NOR2_X1 port map( A1 => n38, A2 => n36, ZN => ab_7_1_port);
   U54 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => ab_7_0_port);
   U55 : NOR2_X1 port map( A1 => n30, A2 => n39, ZN => ab_6_7_port);
   U56 : NOR2_X1 port map( A1 => n33, A2 => n39, ZN => ab_6_6_port);
   U57 : NOR2_X1 port map( A1 => n34, A2 => n39, ZN => ab_6_5_port);
   U58 : NOR2_X1 port map( A1 => n35, A2 => n39, ZN => ab_6_4_port);
   U59 : NOR2_X1 port map( A1 => n31, A2 => n39, ZN => ab_6_3_port);
   U60 : NOR2_X1 port map( A1 => n32, A2 => n39, ZN => ab_6_2_port);
   U61 : NOR2_X1 port map( A1 => n36, A2 => n39, ZN => ab_6_1_port);
   U62 : NOR2_X1 port map( A1 => n37, A2 => n39, ZN => ab_6_0_port);
   U63 : NOR2_X1 port map( A1 => n30, A2 => n40, ZN => ab_5_7_port);
   U64 : NOR2_X1 port map( A1 => n33, A2 => n40, ZN => ab_5_6_port);
   U65 : NOR2_X1 port map( A1 => n34, A2 => n40, ZN => ab_5_5_port);
   U66 : NOR2_X1 port map( A1 => n35, A2 => n40, ZN => ab_5_4_port);
   U67 : NOR2_X1 port map( A1 => n31, A2 => n40, ZN => ab_5_3_port);
   U68 : NOR2_X1 port map( A1 => n32, A2 => n40, ZN => ab_5_2_port);
   U69 : NOR2_X1 port map( A1 => n36, A2 => n40, ZN => ab_5_1_port);
   U70 : NOR2_X1 port map( A1 => n37, A2 => n40, ZN => ab_5_0_port);
   U71 : NOR2_X1 port map( A1 => n30, A2 => n41, ZN => ab_4_7_port);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n41, ZN => ab_4_6_port);
   U73 : NOR2_X1 port map( A1 => n34, A2 => n41, ZN => ab_4_5_port);
   U74 : NOR2_X1 port map( A1 => n35, A2 => n41, ZN => ab_4_4_port);
   U75 : NOR2_X1 port map( A1 => n31, A2 => n41, ZN => ab_4_3_port);
   U76 : NOR2_X1 port map( A1 => n32, A2 => n41, ZN => ab_4_2_port);
   U77 : NOR2_X1 port map( A1 => n36, A2 => n41, ZN => ab_4_1_port);
   U78 : NOR2_X1 port map( A1 => n37, A2 => n41, ZN => ab_4_0_port);
   U79 : NOR2_X1 port map( A1 => n30, A2 => n42, ZN => ab_3_7_port);
   U80 : NOR2_X1 port map( A1 => n33, A2 => n42, ZN => ab_3_6_port);
   U81 : NOR2_X1 port map( A1 => n34, A2 => n42, ZN => ab_3_5_port);
   U82 : NOR2_X1 port map( A1 => n35, A2 => n42, ZN => ab_3_4_port);
   U83 : NOR2_X1 port map( A1 => n31, A2 => n42, ZN => ab_3_3_port);
   U84 : NOR2_X1 port map( A1 => n32, A2 => n42, ZN => ab_3_2_port);
   U85 : NOR2_X1 port map( A1 => n36, A2 => n42, ZN => ab_3_1_port);
   U86 : NOR2_X1 port map( A1 => n37, A2 => n42, ZN => ab_3_0_port);
   U87 : NOR2_X1 port map( A1 => n30, A2 => n43, ZN => ab_2_7_port);
   U88 : NOR2_X1 port map( A1 => n33, A2 => n43, ZN => ab_2_6_port);
   U89 : NOR2_X1 port map( A1 => n34, A2 => n43, ZN => ab_2_5_port);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n43, ZN => ab_2_4_port);
   U91 : NOR2_X1 port map( A1 => n31, A2 => n43, ZN => ab_2_3_port);
   U92 : NOR2_X1 port map( A1 => n32, A2 => n43, ZN => ab_2_2_port);
   U93 : NOR2_X1 port map( A1 => n36, A2 => n43, ZN => ab_2_1_port);
   U94 : NOR2_X1 port map( A1 => n37, A2 => n43, ZN => ab_2_0_port);
   U95 : NOR2_X1 port map( A1 => n30, A2 => n44, ZN => ab_1_7_port);
   U96 : NOR2_X1 port map( A1 => n33, A2 => n44, ZN => ab_1_6_port);
   U97 : NOR2_X1 port map( A1 => n34, A2 => n44, ZN => ab_1_5_port);
   U98 : NOR2_X1 port map( A1 => n35, A2 => n44, ZN => ab_1_4_port);
   U99 : NOR2_X1 port map( A1 => n31, A2 => n44, ZN => ab_1_3_port);
   U100 : NOR2_X1 port map( A1 => n32, A2 => n44, ZN => ab_1_2_port);
   U101 : NOR2_X1 port map( A1 => n36, A2 => n44, ZN => ab_1_1_port);
   U102 : NOR2_X1 port map( A1 => n37, A2 => n44, ZN => ab_1_0_port);
   U103 : NOR2_X1 port map( A1 => n30, A2 => n45, ZN => ab_0_7_port);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n45, ZN => ab_0_6_port);
   U105 : NOR2_X1 port map( A1 => n34, A2 => n45, ZN => ab_0_5_port);
   U106 : NOR2_X1 port map( A1 => n35, A2 => n45, ZN => ab_0_4_port);
   U107 : NOR2_X1 port map( A1 => n31, A2 => n45, ZN => ab_0_3_port);
   U108 : NOR2_X1 port map( A1 => n32, A2 => n45, ZN => ab_0_2_port);
   U109 : NOR2_X1 port map( A1 => n36, A2 => n45, ZN => ab_0_1_port);
   U110 : NOR2_X1 port map( A1 => n37, A2 => n45, ZN => PRODUCT(0));
   n47 <= '0';

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_3_DW01_add_0_DW01_add_2 is

   port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (13 downto 0);  CO : out std_logic);

end shift_pow2_N8_3_DW01_add_0_DW01_add_2;

architecture SYN_cla of shift_pow2_N8_3_DW01_add_0_DW01_add_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, n1, SUM_7_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SUM <= ( SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, SUM_7_port, A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n1);
   U3 : INV_X1 port map( A => n24, ZN => n4);
   U4 : INV_X1 port map( A => n12, ZN => n7);
   U5 : INV_X1 port map( A => n27, ZN => n5);
   U6 : INV_X1 port map( A => n16, ZN => n8);
   U7 : INV_X1 port map( A => n32, ZN => n6);
   U8 : INV_X1 port map( A => n20, ZN => n3);
   U9 : XNOR2_X1 port map( A => B(13), B => n17, ZN => SUM_13_port);
   U10 : AND2_X1 port map( A1 => n16, A2 => n1, ZN => SUM_7_port);
   U11 : XNOR2_X1 port map( A => n9, B => n10, ZN => SUM_9_port);
   U12 : NOR2_X1 port map( A1 => n7, A2 => n11, ZN => n10);
   U13 : XOR2_X1 port map( A => n8, B => n13, Z => SUM_8_port);
   U14 : AND2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U15 : AOI21_X1 port map( B1 => n18, B2 => n3, A => n19, ZN => n17);
   U16 : XOR2_X1 port map( A => n18, B => n21, Z => SUM_12_port);
   U17 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U18 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n19);
   U19 : NOR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n20);
   U20 : OAI211_X1 port map( C1 => n22, C2 => n23, A => n24, B => n25, ZN => 
                           n18);
   U21 : OR4_X1 port map( A1 => n26, A2 => n27, A3 => n23, A4 => n11, ZN => n25
                           );
   U22 : AOI21_X1 port map( B1 => n5, B2 => n28, A => n6, ZN => n22);
   U23 : OAI21_X1 port map( B1 => n11, B2 => n15, A => n12, ZN => n28);
   U24 : XNOR2_X1 port map( A => n29, B => n30, ZN => SUM_11_port);
   U25 : NOR2_X1 port map( A1 => n23, A2 => n4, ZN => n30);
   U26 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n24);
   U27 : NOR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n23);
   U28 : AOI21_X1 port map( B1 => n31, B2 => n5, A => n6, ZN => n29);
   U29 : XNOR2_X1 port map( A => n33, B => n31, ZN => SUM_10_port);
   U30 : OAI21_X1 port map( B1 => n11, B2 => n9, A => n12, ZN => n31);
   U31 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n12);
   U32 : AND2_X1 port map( A1 => n26, A2 => n15, ZN => n9);
   U33 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n15);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n14, ZN => n26);
   U35 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n14);
   U36 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n16);
   U37 : NOR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n11);
   U38 : NAND2_X1 port map( A1 => n32, A2 => n5, ZN => n33);
   U39 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n27);
   U40 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n32);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_3_DW02_mult_0_DW02_mult_2 is

   port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  PRODUCT 
         : out std_logic_vector (15 downto 0));

end shift_pow2_N8_3_DW02_mult_0_DW02_mult_2;

architecture SYN_csa of shift_pow2_N8_3_DW02_mult_0_DW02_mult_2 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component shift_pow2_N8_3_DW01_add_0_DW01_add_2
      port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (13 downto 0);  CO : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, ab_7_4_port, 
      ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_7_port, ab_3_6_port, 
      ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, 
      ab_3_0_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, ab_2_4_port, 
      ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, ab_1_7_port, 
      ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_2_port, 
      ab_1_1_port, ab_1_0_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, 
      SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, SUMB_7_0_port, SUMB_6_6_port
      , SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, 
      SUMB_6_1_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_6_port, SUMB_4_5_port, 
      SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_6_port
      , SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, 
      SUMB_3_1_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n_1071 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => 
                           SUMB_7_0_port);
   S4_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S4_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S4_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S4_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S4_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S5_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           ab_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S3_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           ab_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S3_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           ab_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S3_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           ab_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S3_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           ab_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n7, CI => n13, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n6, CI => n12, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n5, CI => n11, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n4, CI => n10, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n3, CI => n14, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n2, CI => n9, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S3_2_6 : FA_X1 port map( A => ab_2_6_port, B => n8, CI => ab_1_7_port, CO =>
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   FS_1 : shift_pow2_N8_3_DW01_add_0_DW01_add_2 port map( A(13) => n46, A(12) 
                           => n17, A(11) => n20, A(10) => n19, A(9) => n22, 
                           A(8) => n27, A(7) => n21, A(6) => n18, A(5) => 
                           SUMB_7_0_port, A(4) => A1_4_port, A(3) => A1_3_port,
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(13) => n15, B(12) => n28, B(11) => n25,
                           B(10) => n24, B(9) => n26, B(8) => n29, B(7) => n23,
                           B(6) => n46, B(5) => n47, B(4) => n47, B(3) => n47, 
                           B(2) => n47, B(1) => n47, B(0) => X_Logic0_port, CI 
                           => X_Logic0_port, SUM(13) => PRODUCT(15), SUM(12) =>
                           PRODUCT(14), SUM(11) => PRODUCT(13), SUM(10) => 
                           PRODUCT(12), SUM(9) => PRODUCT(11), SUM(8) => 
                           PRODUCT(10), SUM(7) => PRODUCT(9), SUM(6) => 
                           PRODUCT(8), SUM(5) => PRODUCT(7), SUM(4) => 
                           PRODUCT(6), SUM(3) => PRODUCT(5), SUM(2) => 
                           PRODUCT(4), SUM(1) => PRODUCT(3), SUM(0) => 
                           PRODUCT(2), CO => n_1071);
   U2 : INV_X1 port map( A => B(4), ZN => n35);
   U3 : INV_X1 port map( A => B(5), ZN => n34);
   U4 : INV_X1 port map( A => B(6), ZN => n33);
   U5 : INV_X1 port map( A => B(7), ZN => n30);
   U6 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n2);
   U7 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n3);
   U8 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n4);
   U9 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n5);
   U10 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n6);
   U11 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n7);
   U12 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n8);
   U13 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n9);
   U14 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n10);
   U15 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n11);
   U16 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n12);
   U17 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n13);
   U18 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n14);
   U19 : AND2_X1 port map( A1 => CARRYB_7_6_port, A2 => ab_7_7_port, ZN => n15)
                           ;
   U20 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U21 : XOR2_X1 port map( A => CARRYB_7_6_port, B => ab_7_7_port, Z => n17);
   U22 : XOR2_X1 port map( A => CARRYB_7_0_port, B => SUMB_7_1_port, Z => n18);
   U23 : XOR2_X1 port map( A => CARRYB_7_4_port, B => SUMB_7_5_port, Z => n19);
   U24 : XOR2_X1 port map( A => CARRYB_7_5_port, B => SUMB_7_6_port, Z => n20);
   U25 : XOR2_X1 port map( A => CARRYB_7_1_port, B => SUMB_7_2_port, Z => n21);
   U26 : XOR2_X1 port map( A => CARRYB_7_3_port, B => SUMB_7_4_port, Z => n22);
   U27 : AND2_X1 port map( A1 => CARRYB_7_0_port, A2 => SUMB_7_1_port, ZN => 
                           n23);
   U28 : AND2_X1 port map( A1 => CARRYB_7_3_port, A2 => SUMB_7_4_port, ZN => 
                           n24);
   U29 : AND2_X1 port map( A1 => CARRYB_7_4_port, A2 => SUMB_7_5_port, ZN => 
                           n25);
   U30 : AND2_X1 port map( A1 => CARRYB_7_2_port, A2 => SUMB_7_3_port, ZN => 
                           n26);
   U31 : XOR2_X1 port map( A => CARRYB_7_2_port, B => SUMB_7_3_port, Z => n27);
   U32 : AND2_X1 port map( A1 => CARRYB_7_5_port, A2 => SUMB_7_6_port, ZN => 
                           n28);
   U33 : AND2_X1 port map( A1 => CARRYB_7_1_port, A2 => SUMB_7_2_port, ZN => 
                           n29);
   U34 : INV_X1 port map( A => B(2), ZN => n32);
   U35 : INV_X1 port map( A => B(1), ZN => n36);
   U36 : INV_X1 port map( A => B(0), ZN => n37);
   U37 : INV_X1 port map( A => B(3), ZN => n31);
   U38 : INV_X1 port map( A => A(7), ZN => n38);
   U39 : INV_X1 port map( A => A(0), ZN => n45);
   U40 : INV_X1 port map( A => A(1), ZN => n44);
   U41 : INV_X1 port map( A => A(2), ZN => n43);
   U42 : INV_X1 port map( A => A(3), ZN => n42);
   U43 : INV_X1 port map( A => A(4), ZN => n41);
   U44 : INV_X1 port map( A => A(5), ZN => n40);
   U45 : INV_X1 port map( A => A(6), ZN => n39);
   n46 <= '0';
   U47 : NOR2_X1 port map( A1 => n38, A2 => n30, ZN => ab_7_7_port);
   U48 : NOR2_X1 port map( A1 => n38, A2 => n33, ZN => ab_7_6_port);
   U49 : NOR2_X1 port map( A1 => n38, A2 => n34, ZN => ab_7_5_port);
   U50 : NOR2_X1 port map( A1 => n38, A2 => n35, ZN => ab_7_4_port);
   U51 : NOR2_X1 port map( A1 => n38, A2 => n31, ZN => ab_7_3_port);
   U52 : NOR2_X1 port map( A1 => n38, A2 => n32, ZN => ab_7_2_port);
   U53 : NOR2_X1 port map( A1 => n38, A2 => n36, ZN => ab_7_1_port);
   U54 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => ab_7_0_port);
   U55 : NOR2_X1 port map( A1 => n30, A2 => n39, ZN => ab_6_7_port);
   U56 : NOR2_X1 port map( A1 => n33, A2 => n39, ZN => ab_6_6_port);
   U57 : NOR2_X1 port map( A1 => n34, A2 => n39, ZN => ab_6_5_port);
   U58 : NOR2_X1 port map( A1 => n35, A2 => n39, ZN => ab_6_4_port);
   U59 : NOR2_X1 port map( A1 => n31, A2 => n39, ZN => ab_6_3_port);
   U60 : NOR2_X1 port map( A1 => n32, A2 => n39, ZN => ab_6_2_port);
   U61 : NOR2_X1 port map( A1 => n36, A2 => n39, ZN => ab_6_1_port);
   U62 : NOR2_X1 port map( A1 => n37, A2 => n39, ZN => ab_6_0_port);
   U63 : NOR2_X1 port map( A1 => n30, A2 => n40, ZN => ab_5_7_port);
   U64 : NOR2_X1 port map( A1 => n33, A2 => n40, ZN => ab_5_6_port);
   U65 : NOR2_X1 port map( A1 => n34, A2 => n40, ZN => ab_5_5_port);
   U66 : NOR2_X1 port map( A1 => n35, A2 => n40, ZN => ab_5_4_port);
   U67 : NOR2_X1 port map( A1 => n31, A2 => n40, ZN => ab_5_3_port);
   U68 : NOR2_X1 port map( A1 => n32, A2 => n40, ZN => ab_5_2_port);
   U69 : NOR2_X1 port map( A1 => n36, A2 => n40, ZN => ab_5_1_port);
   U70 : NOR2_X1 port map( A1 => n37, A2 => n40, ZN => ab_5_0_port);
   U71 : NOR2_X1 port map( A1 => n30, A2 => n41, ZN => ab_4_7_port);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n41, ZN => ab_4_6_port);
   U73 : NOR2_X1 port map( A1 => n34, A2 => n41, ZN => ab_4_5_port);
   U74 : NOR2_X1 port map( A1 => n35, A2 => n41, ZN => ab_4_4_port);
   U75 : NOR2_X1 port map( A1 => n31, A2 => n41, ZN => ab_4_3_port);
   U76 : NOR2_X1 port map( A1 => n32, A2 => n41, ZN => ab_4_2_port);
   U77 : NOR2_X1 port map( A1 => n36, A2 => n41, ZN => ab_4_1_port);
   U78 : NOR2_X1 port map( A1 => n37, A2 => n41, ZN => ab_4_0_port);
   U79 : NOR2_X1 port map( A1 => n30, A2 => n42, ZN => ab_3_7_port);
   U80 : NOR2_X1 port map( A1 => n33, A2 => n42, ZN => ab_3_6_port);
   U81 : NOR2_X1 port map( A1 => n34, A2 => n42, ZN => ab_3_5_port);
   U82 : NOR2_X1 port map( A1 => n35, A2 => n42, ZN => ab_3_4_port);
   U83 : NOR2_X1 port map( A1 => n31, A2 => n42, ZN => ab_3_3_port);
   U84 : NOR2_X1 port map( A1 => n32, A2 => n42, ZN => ab_3_2_port);
   U85 : NOR2_X1 port map( A1 => n36, A2 => n42, ZN => ab_3_1_port);
   U86 : NOR2_X1 port map( A1 => n37, A2 => n42, ZN => ab_3_0_port);
   U87 : NOR2_X1 port map( A1 => n30, A2 => n43, ZN => ab_2_7_port);
   U88 : NOR2_X1 port map( A1 => n33, A2 => n43, ZN => ab_2_6_port);
   U89 : NOR2_X1 port map( A1 => n34, A2 => n43, ZN => ab_2_5_port);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n43, ZN => ab_2_4_port);
   U91 : NOR2_X1 port map( A1 => n31, A2 => n43, ZN => ab_2_3_port);
   U92 : NOR2_X1 port map( A1 => n32, A2 => n43, ZN => ab_2_2_port);
   U93 : NOR2_X1 port map( A1 => n36, A2 => n43, ZN => ab_2_1_port);
   U94 : NOR2_X1 port map( A1 => n37, A2 => n43, ZN => ab_2_0_port);
   U95 : NOR2_X1 port map( A1 => n30, A2 => n44, ZN => ab_1_7_port);
   U96 : NOR2_X1 port map( A1 => n33, A2 => n44, ZN => ab_1_6_port);
   U97 : NOR2_X1 port map( A1 => n34, A2 => n44, ZN => ab_1_5_port);
   U98 : NOR2_X1 port map( A1 => n35, A2 => n44, ZN => ab_1_4_port);
   U99 : NOR2_X1 port map( A1 => n31, A2 => n44, ZN => ab_1_3_port);
   U100 : NOR2_X1 port map( A1 => n32, A2 => n44, ZN => ab_1_2_port);
   U101 : NOR2_X1 port map( A1 => n36, A2 => n44, ZN => ab_1_1_port);
   U102 : NOR2_X1 port map( A1 => n37, A2 => n44, ZN => ab_1_0_port);
   U103 : NOR2_X1 port map( A1 => n30, A2 => n45, ZN => ab_0_7_port);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n45, ZN => ab_0_6_port);
   U105 : NOR2_X1 port map( A1 => n34, A2 => n45, ZN => ab_0_5_port);
   U106 : NOR2_X1 port map( A1 => n35, A2 => n45, ZN => ab_0_4_port);
   U107 : NOR2_X1 port map( A1 => n31, A2 => n45, ZN => ab_0_3_port);
   U108 : NOR2_X1 port map( A1 => n32, A2 => n45, ZN => ab_0_2_port);
   U109 : NOR2_X1 port map( A1 => n36, A2 => n45, ZN => ab_0_1_port);
   U110 : NOR2_X1 port map( A1 => n37, A2 => n45, ZN => PRODUCT(0));
   n47 <= '0';

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_2_DW01_add_0_DW01_add_1 is

   port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (13 downto 0);  CO : out std_logic);

end shift_pow2_N8_2_DW01_add_0_DW01_add_1;

architecture SYN_cla of shift_pow2_N8_2_DW01_add_0_DW01_add_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, n1, SUM_7_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SUM <= ( SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, SUM_7_port, A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n1);
   U3 : INV_X1 port map( A => n24, ZN => n4);
   U4 : INV_X1 port map( A => n12, ZN => n7);
   U5 : INV_X1 port map( A => n27, ZN => n5);
   U6 : INV_X1 port map( A => n16, ZN => n8);
   U7 : INV_X1 port map( A => n32, ZN => n6);
   U8 : INV_X1 port map( A => n20, ZN => n3);
   U9 : XNOR2_X1 port map( A => B(13), B => n17, ZN => SUM_13_port);
   U10 : AND2_X1 port map( A1 => n16, A2 => n1, ZN => SUM_7_port);
   U11 : XNOR2_X1 port map( A => n9, B => n10, ZN => SUM_9_port);
   U12 : NOR2_X1 port map( A1 => n7, A2 => n11, ZN => n10);
   U13 : XOR2_X1 port map( A => n8, B => n13, Z => SUM_8_port);
   U14 : AND2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U15 : AOI21_X1 port map( B1 => n18, B2 => n3, A => n19, ZN => n17);
   U16 : XOR2_X1 port map( A => n18, B => n21, Z => SUM_12_port);
   U17 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U18 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n19);
   U19 : NOR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n20);
   U20 : OAI211_X1 port map( C1 => n22, C2 => n23, A => n24, B => n25, ZN => 
                           n18);
   U21 : OR4_X1 port map( A1 => n26, A2 => n27, A3 => n23, A4 => n11, ZN => n25
                           );
   U22 : AOI21_X1 port map( B1 => n5, B2 => n28, A => n6, ZN => n22);
   U23 : OAI21_X1 port map( B1 => n11, B2 => n15, A => n12, ZN => n28);
   U24 : XNOR2_X1 port map( A => n29, B => n30, ZN => SUM_11_port);
   U25 : NOR2_X1 port map( A1 => n23, A2 => n4, ZN => n30);
   U26 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n24);
   U27 : NOR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n23);
   U28 : AOI21_X1 port map( B1 => n31, B2 => n5, A => n6, ZN => n29);
   U29 : XNOR2_X1 port map( A => n33, B => n31, ZN => SUM_10_port);
   U30 : OAI21_X1 port map( B1 => n11, B2 => n9, A => n12, ZN => n31);
   U31 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n12);
   U32 : AND2_X1 port map( A1 => n26, A2 => n15, ZN => n9);
   U33 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n15);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n14, ZN => n26);
   U35 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n14);
   U36 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n16);
   U37 : NOR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n11);
   U38 : NAND2_X1 port map( A1 => n32, A2 => n5, ZN => n33);
   U39 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n27);
   U40 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n32);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_2_DW02_mult_0_DW02_mult_1 is

   port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  PRODUCT 
         : out std_logic_vector (15 downto 0));

end shift_pow2_N8_2_DW02_mult_0_DW02_mult_1;

architecture SYN_csa of shift_pow2_N8_2_DW02_mult_0_DW02_mult_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component shift_pow2_N8_2_DW01_add_0_DW01_add_1
      port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (13 downto 0);  CO : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, ab_7_4_port, 
      ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_7_port, ab_3_6_port, 
      ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, 
      ab_3_0_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, ab_2_4_port, 
      ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, ab_1_7_port, 
      ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_2_port, 
      ab_1_1_port, ab_1_0_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, 
      SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, SUMB_7_0_port, SUMB_6_6_port
      , SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, 
      SUMB_6_1_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_6_port, SUMB_4_5_port, 
      SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_6_port
      , SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, 
      SUMB_3_1_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n_1083 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => 
                           SUMB_7_0_port);
   S4_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S4_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S4_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S4_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S4_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S5_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           ab_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S3_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           ab_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S3_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           ab_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S3_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           ab_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S3_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           ab_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n7, CI => n13, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n6, CI => n12, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n5, CI => n11, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n4, CI => n10, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n3, CI => n9, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n2, CI => n14, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S3_2_6 : FA_X1 port map( A => ab_2_6_port, B => n8, CI => ab_1_7_port, CO =>
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   FS_1 : shift_pow2_N8_2_DW01_add_0_DW01_add_1 port map( A(13) => n46, A(12) 
                           => n18, A(11) => n19, A(10) => n21, A(9) => n22, 
                           A(8) => n27, A(7) => n20, A(6) => n17, A(5) => 
                           SUMB_7_0_port, A(4) => A1_4_port, A(3) => A1_3_port,
                           A(2) => A1_2_port, A(1) => A1_1_port, A(0) => 
                           A1_0_port, B(13) => n15, B(12) => n28, B(11) => n25,
                           B(10) => n24, B(9) => n26, B(8) => n29, B(7) => n23,
                           B(6) => n46, B(5) => n47, B(4) => n47, B(3) => n47, 
                           B(2) => n47, B(1) => n47, B(0) => X_Logic0_port, CI 
                           => X_Logic0_port, SUM(13) => PRODUCT(15), SUM(12) =>
                           PRODUCT(14), SUM(11) => PRODUCT(13), SUM(10) => 
                           PRODUCT(12), SUM(9) => PRODUCT(11), SUM(8) => 
                           PRODUCT(10), SUM(7) => PRODUCT(9), SUM(6) => 
                           PRODUCT(8), SUM(5) => PRODUCT(7), SUM(4) => 
                           PRODUCT(6), SUM(3) => PRODUCT(5), SUM(2) => 
                           PRODUCT(4), SUM(1) => PRODUCT(3), SUM(0) => 
                           PRODUCT(2), CO => n_1083);
   U2 : INV_X1 port map( A => B(4), ZN => n35);
   U3 : INV_X1 port map( A => B(5), ZN => n34);
   U4 : INV_X1 port map( A => B(6), ZN => n33);
   U5 : INV_X1 port map( A => B(7), ZN => n30);
   U6 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n2);
   U7 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n3);
   U8 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n4);
   U9 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n5);
   U10 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n6);
   U11 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n7);
   U12 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n8);
   U13 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n9);
   U14 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n10);
   U15 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n11);
   U16 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n12);
   U17 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n13);
   U18 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n14);
   U19 : AND2_X1 port map( A1 => CARRYB_7_6_port, A2 => ab_7_7_port, ZN => n15)
                           ;
   U20 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U21 : XOR2_X1 port map( A => CARRYB_7_0_port, B => SUMB_7_1_port, Z => n17);
   U22 : XOR2_X1 port map( A => CARRYB_7_6_port, B => ab_7_7_port, Z => n18);
   U23 : XOR2_X1 port map( A => CARRYB_7_5_port, B => SUMB_7_6_port, Z => n19);
   U24 : XOR2_X1 port map( A => CARRYB_7_1_port, B => SUMB_7_2_port, Z => n20);
   U25 : XOR2_X1 port map( A => CARRYB_7_4_port, B => SUMB_7_5_port, Z => n21);
   U26 : XOR2_X1 port map( A => CARRYB_7_3_port, B => SUMB_7_4_port, Z => n22);
   U27 : AND2_X1 port map( A1 => CARRYB_7_0_port, A2 => SUMB_7_1_port, ZN => 
                           n23);
   U28 : AND2_X1 port map( A1 => CARRYB_7_3_port, A2 => SUMB_7_4_port, ZN => 
                           n24);
   U29 : AND2_X1 port map( A1 => CARRYB_7_4_port, A2 => SUMB_7_5_port, ZN => 
                           n25);
   U30 : AND2_X1 port map( A1 => CARRYB_7_2_port, A2 => SUMB_7_3_port, ZN => 
                           n26);
   U31 : XOR2_X1 port map( A => CARRYB_7_2_port, B => SUMB_7_3_port, Z => n27);
   U32 : AND2_X1 port map( A1 => CARRYB_7_5_port, A2 => SUMB_7_6_port, ZN => 
                           n28);
   U33 : AND2_X1 port map( A1 => CARRYB_7_1_port, A2 => SUMB_7_2_port, ZN => 
                           n29);
   U34 : INV_X1 port map( A => B(2), ZN => n32);
   U35 : INV_X1 port map( A => B(1), ZN => n36);
   U36 : INV_X1 port map( A => B(3), ZN => n31);
   U37 : INV_X1 port map( A => B(0), ZN => n37);
   U38 : INV_X1 port map( A => A(7), ZN => n38);
   U39 : INV_X1 port map( A => A(0), ZN => n45);
   U40 : INV_X1 port map( A => A(1), ZN => n44);
   U41 : INV_X1 port map( A => A(3), ZN => n42);
   U42 : INV_X1 port map( A => A(4), ZN => n41);
   U43 : INV_X1 port map( A => A(5), ZN => n40);
   U44 : INV_X1 port map( A => A(6), ZN => n39);
   U45 : INV_X1 port map( A => A(2), ZN => n43);
   n46 <= '0';
   U47 : NOR2_X1 port map( A1 => n38, A2 => n30, ZN => ab_7_7_port);
   U48 : NOR2_X1 port map( A1 => n38, A2 => n33, ZN => ab_7_6_port);
   U49 : NOR2_X1 port map( A1 => n38, A2 => n34, ZN => ab_7_5_port);
   U50 : NOR2_X1 port map( A1 => n38, A2 => n35, ZN => ab_7_4_port);
   U51 : NOR2_X1 port map( A1 => n38, A2 => n31, ZN => ab_7_3_port);
   U52 : NOR2_X1 port map( A1 => n38, A2 => n32, ZN => ab_7_2_port);
   U53 : NOR2_X1 port map( A1 => n38, A2 => n36, ZN => ab_7_1_port);
   U54 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => ab_7_0_port);
   U55 : NOR2_X1 port map( A1 => n30, A2 => n39, ZN => ab_6_7_port);
   U56 : NOR2_X1 port map( A1 => n33, A2 => n39, ZN => ab_6_6_port);
   U57 : NOR2_X1 port map( A1 => n34, A2 => n39, ZN => ab_6_5_port);
   U58 : NOR2_X1 port map( A1 => n35, A2 => n39, ZN => ab_6_4_port);
   U59 : NOR2_X1 port map( A1 => n31, A2 => n39, ZN => ab_6_3_port);
   U60 : NOR2_X1 port map( A1 => n32, A2 => n39, ZN => ab_6_2_port);
   U61 : NOR2_X1 port map( A1 => n36, A2 => n39, ZN => ab_6_1_port);
   U62 : NOR2_X1 port map( A1 => n37, A2 => n39, ZN => ab_6_0_port);
   U63 : NOR2_X1 port map( A1 => n30, A2 => n40, ZN => ab_5_7_port);
   U64 : NOR2_X1 port map( A1 => n33, A2 => n40, ZN => ab_5_6_port);
   U65 : NOR2_X1 port map( A1 => n34, A2 => n40, ZN => ab_5_5_port);
   U66 : NOR2_X1 port map( A1 => n35, A2 => n40, ZN => ab_5_4_port);
   U67 : NOR2_X1 port map( A1 => n31, A2 => n40, ZN => ab_5_3_port);
   U68 : NOR2_X1 port map( A1 => n32, A2 => n40, ZN => ab_5_2_port);
   U69 : NOR2_X1 port map( A1 => n36, A2 => n40, ZN => ab_5_1_port);
   U70 : NOR2_X1 port map( A1 => n37, A2 => n40, ZN => ab_5_0_port);
   U71 : NOR2_X1 port map( A1 => n30, A2 => n41, ZN => ab_4_7_port);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n41, ZN => ab_4_6_port);
   U73 : NOR2_X1 port map( A1 => n34, A2 => n41, ZN => ab_4_5_port);
   U74 : NOR2_X1 port map( A1 => n35, A2 => n41, ZN => ab_4_4_port);
   U75 : NOR2_X1 port map( A1 => n31, A2 => n41, ZN => ab_4_3_port);
   U76 : NOR2_X1 port map( A1 => n32, A2 => n41, ZN => ab_4_2_port);
   U77 : NOR2_X1 port map( A1 => n36, A2 => n41, ZN => ab_4_1_port);
   U78 : NOR2_X1 port map( A1 => n37, A2 => n41, ZN => ab_4_0_port);
   U79 : NOR2_X1 port map( A1 => n30, A2 => n42, ZN => ab_3_7_port);
   U80 : NOR2_X1 port map( A1 => n33, A2 => n42, ZN => ab_3_6_port);
   U81 : NOR2_X1 port map( A1 => n34, A2 => n42, ZN => ab_3_5_port);
   U82 : NOR2_X1 port map( A1 => n35, A2 => n42, ZN => ab_3_4_port);
   U83 : NOR2_X1 port map( A1 => n31, A2 => n42, ZN => ab_3_3_port);
   U84 : NOR2_X1 port map( A1 => n32, A2 => n42, ZN => ab_3_2_port);
   U85 : NOR2_X1 port map( A1 => n36, A2 => n42, ZN => ab_3_1_port);
   U86 : NOR2_X1 port map( A1 => n37, A2 => n42, ZN => ab_3_0_port);
   U87 : NOR2_X1 port map( A1 => n30, A2 => n43, ZN => ab_2_7_port);
   U88 : NOR2_X1 port map( A1 => n33, A2 => n43, ZN => ab_2_6_port);
   U89 : NOR2_X1 port map( A1 => n34, A2 => n43, ZN => ab_2_5_port);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n43, ZN => ab_2_4_port);
   U91 : NOR2_X1 port map( A1 => n31, A2 => n43, ZN => ab_2_3_port);
   U92 : NOR2_X1 port map( A1 => n32, A2 => n43, ZN => ab_2_2_port);
   U93 : NOR2_X1 port map( A1 => n36, A2 => n43, ZN => ab_2_1_port);
   U94 : NOR2_X1 port map( A1 => n37, A2 => n43, ZN => ab_2_0_port);
   U95 : NOR2_X1 port map( A1 => n30, A2 => n44, ZN => ab_1_7_port);
   U96 : NOR2_X1 port map( A1 => n33, A2 => n44, ZN => ab_1_6_port);
   U97 : NOR2_X1 port map( A1 => n34, A2 => n44, ZN => ab_1_5_port);
   U98 : NOR2_X1 port map( A1 => n35, A2 => n44, ZN => ab_1_4_port);
   U99 : NOR2_X1 port map( A1 => n31, A2 => n44, ZN => ab_1_3_port);
   U100 : NOR2_X1 port map( A1 => n32, A2 => n44, ZN => ab_1_2_port);
   U101 : NOR2_X1 port map( A1 => n36, A2 => n44, ZN => ab_1_1_port);
   U102 : NOR2_X1 port map( A1 => n37, A2 => n44, ZN => ab_1_0_port);
   U103 : NOR2_X1 port map( A1 => n30, A2 => n45, ZN => ab_0_7_port);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n45, ZN => ab_0_6_port);
   U105 : NOR2_X1 port map( A1 => n34, A2 => n45, ZN => ab_0_5_port);
   U106 : NOR2_X1 port map( A1 => n35, A2 => n45, ZN => ab_0_4_port);
   U107 : NOR2_X1 port map( A1 => n31, A2 => n45, ZN => ab_0_3_port);
   U108 : NOR2_X1 port map( A1 => n32, A2 => n45, ZN => ab_0_2_port);
   U109 : NOR2_X1 port map( A1 => n36, A2 => n45, ZN => ab_0_1_port);
   U110 : NOR2_X1 port map( A1 => n37, A2 => n45, ZN => PRODUCT(0));
   n47 <= '0';

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_1_DW01_add_0 is

   port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (13 downto 0);  CO : out std_logic);

end shift_pow2_N8_1_DW01_add_0;

architecture SYN_cla of shift_pow2_N8_1_DW01_add_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, n1, SUM_7_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33 : std_logic;

begin
   SUM <= ( SUM_13_port, SUM_12_port, SUM_11_port, SUM_10_port, SUM_9_port, 
      SUM_8_port, SUM_7_port, A(6), A(5), A(4), A(3), A(2), A(1), A(0) );
   
   U2 : OR2_X1 port map( A1 => B(7), A2 => A(7), ZN => n1);
   U3 : INV_X1 port map( A => n24, ZN => n4);
   U4 : INV_X1 port map( A => n12, ZN => n7);
   U5 : INV_X1 port map( A => n27, ZN => n5);
   U6 : INV_X1 port map( A => n16, ZN => n8);
   U7 : INV_X1 port map( A => n32, ZN => n6);
   U8 : INV_X1 port map( A => n20, ZN => n3);
   U9 : XNOR2_X1 port map( A => B(13), B => n17, ZN => SUM_13_port);
   U10 : AND2_X1 port map( A1 => n16, A2 => n1, ZN => SUM_7_port);
   U11 : XNOR2_X1 port map( A => n9, B => n10, ZN => SUM_9_port);
   U12 : NOR2_X1 port map( A1 => n7, A2 => n11, ZN => n10);
   U13 : XOR2_X1 port map( A => n8, B => n13, Z => SUM_8_port);
   U14 : AND2_X1 port map( A1 => n14, A2 => n15, ZN => n13);
   U15 : AOI21_X1 port map( B1 => n18, B2 => n3, A => n19, ZN => n17);
   U16 : XOR2_X1 port map( A => n18, B => n21, Z => SUM_12_port);
   U17 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U18 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n19);
   U19 : NOR2_X1 port map( A1 => B(12), A2 => A(12), ZN => n20);
   U20 : OAI211_X1 port map( C1 => n22, C2 => n23, A => n24, B => n25, ZN => 
                           n18);
   U21 : OR4_X1 port map( A1 => n26, A2 => n27, A3 => n23, A4 => n11, ZN => n25
                           );
   U22 : AOI21_X1 port map( B1 => n5, B2 => n28, A => n6, ZN => n22);
   U23 : OAI21_X1 port map( B1 => n11, B2 => n15, A => n12, ZN => n28);
   U24 : XNOR2_X1 port map( A => n29, B => n30, ZN => SUM_11_port);
   U25 : NOR2_X1 port map( A1 => n23, A2 => n4, ZN => n30);
   U26 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n24);
   U27 : NOR2_X1 port map( A1 => B(11), A2 => A(11), ZN => n23);
   U28 : AOI21_X1 port map( B1 => n31, B2 => n5, A => n6, ZN => n29);
   U29 : XNOR2_X1 port map( A => n33, B => n31, ZN => SUM_10_port);
   U30 : OAI21_X1 port map( B1 => n11, B2 => n9, A => n12, ZN => n31);
   U31 : NAND2_X1 port map( A1 => B(9), A2 => A(9), ZN => n12);
   U32 : AND2_X1 port map( A1 => n26, A2 => n15, ZN => n9);
   U33 : NAND2_X1 port map( A1 => B(8), A2 => A(8), ZN => n15);
   U34 : NAND2_X1 port map( A1 => n8, A2 => n14, ZN => n26);
   U35 : OR2_X1 port map( A1 => B(8), A2 => A(8), ZN => n14);
   U36 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n16);
   U37 : NOR2_X1 port map( A1 => B(9), A2 => A(9), ZN => n11);
   U38 : NAND2_X1 port map( A1 => n32, A2 => n5, ZN => n33);
   U39 : NOR2_X1 port map( A1 => B(10), A2 => A(10), ZN => n27);
   U40 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n32);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_1_DW02_mult_0 is

   port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  PRODUCT 
         : out std_logic_vector (15 downto 0));

end shift_pow2_N8_1_DW02_mult_0;

architecture SYN_csa of shift_pow2_N8_1_DW02_mult_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component shift_pow2_N8_1_DW01_add_0
      port( A, B : in std_logic_vector (13 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (13 downto 0);  CO : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal X_Logic0_port, ab_7_7_port, ab_7_6_port, ab_7_5_port, ab_7_4_port, 
      ab_7_3_port, ab_7_2_port, ab_7_1_port, ab_7_0_port, ab_6_7_port, 
      ab_6_6_port, ab_6_5_port, ab_6_4_port, ab_6_3_port, ab_6_2_port, 
      ab_6_1_port, ab_6_0_port, ab_5_7_port, ab_5_6_port, ab_5_5_port, 
      ab_5_4_port, ab_5_3_port, ab_5_2_port, ab_5_1_port, ab_5_0_port, 
      ab_4_7_port, ab_4_6_port, ab_4_5_port, ab_4_4_port, ab_4_3_port, 
      ab_4_2_port, ab_4_1_port, ab_4_0_port, ab_3_7_port, ab_3_6_port, 
      ab_3_5_port, ab_3_4_port, ab_3_3_port, ab_3_2_port, ab_3_1_port, 
      ab_3_0_port, ab_2_7_port, ab_2_6_port, ab_2_5_port, ab_2_4_port, 
      ab_2_3_port, ab_2_2_port, ab_2_1_port, ab_2_0_port, ab_1_7_port, 
      ab_1_6_port, ab_1_5_port, ab_1_4_port, ab_1_3_port, ab_1_2_port, 
      ab_1_1_port, ab_1_0_port, ab_0_7_port, ab_0_6_port, ab_0_5_port, 
      ab_0_4_port, ab_0_3_port, ab_0_2_port, ab_0_1_port, CARRYB_7_6_port, 
      CARRYB_7_5_port, CARRYB_7_4_port, CARRYB_7_3_port, CARRYB_7_2_port, 
      CARRYB_7_1_port, CARRYB_7_0_port, CARRYB_6_6_port, CARRYB_6_5_port, 
      CARRYB_6_4_port, CARRYB_6_3_port, CARRYB_6_2_port, CARRYB_6_1_port, 
      CARRYB_6_0_port, CARRYB_5_6_port, CARRYB_5_5_port, CARRYB_5_4_port, 
      CARRYB_5_3_port, CARRYB_5_2_port, CARRYB_5_1_port, CARRYB_5_0_port, 
      CARRYB_4_6_port, CARRYB_4_5_port, CARRYB_4_4_port, CARRYB_4_3_port, 
      CARRYB_4_2_port, CARRYB_4_1_port, CARRYB_4_0_port, CARRYB_3_6_port, 
      CARRYB_3_5_port, CARRYB_3_4_port, CARRYB_3_3_port, CARRYB_3_2_port, 
      CARRYB_3_1_port, CARRYB_3_0_port, CARRYB_2_6_port, CARRYB_2_5_port, 
      CARRYB_2_4_port, CARRYB_2_3_port, CARRYB_2_2_port, CARRYB_2_1_port, 
      CARRYB_2_0_port, SUMB_7_6_port, SUMB_7_5_port, SUMB_7_4_port, 
      SUMB_7_3_port, SUMB_7_2_port, SUMB_7_1_port, SUMB_7_0_port, SUMB_6_6_port
      , SUMB_6_5_port, SUMB_6_4_port, SUMB_6_3_port, SUMB_6_2_port, 
      SUMB_6_1_port, SUMB_5_6_port, SUMB_5_5_port, SUMB_5_4_port, SUMB_5_3_port
      , SUMB_5_2_port, SUMB_5_1_port, SUMB_4_6_port, SUMB_4_5_port, 
      SUMB_4_4_port, SUMB_4_3_port, SUMB_4_2_port, SUMB_4_1_port, SUMB_3_6_port
      , SUMB_3_5_port, SUMB_3_4_port, SUMB_3_3_port, SUMB_3_2_port, 
      SUMB_3_1_port, SUMB_2_6_port, SUMB_2_5_port, SUMB_2_4_port, SUMB_2_3_port
      , SUMB_2_2_port, SUMB_2_1_port, A1_4_port, A1_3_port, A1_2_port, 
      A1_1_port, A1_0_port, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n_1095 : std_logic;

begin
   
   X_Logic0_port <= '0';
   S4_0 : FA_X1 port map( A => ab_7_0_port, B => CARRYB_6_0_port, CI => 
                           SUMB_6_1_port, CO => CARRYB_7_0_port, S => 
                           SUMB_7_0_port);
   S4_1 : FA_X1 port map( A => ab_7_1_port, B => CARRYB_6_1_port, CI => 
                           SUMB_6_2_port, CO => CARRYB_7_1_port, S => 
                           SUMB_7_1_port);
   S4_2 : FA_X1 port map( A => ab_7_2_port, B => CARRYB_6_2_port, CI => 
                           SUMB_6_3_port, CO => CARRYB_7_2_port, S => 
                           SUMB_7_2_port);
   S4_3 : FA_X1 port map( A => ab_7_3_port, B => CARRYB_6_3_port, CI => 
                           SUMB_6_4_port, CO => CARRYB_7_3_port, S => 
                           SUMB_7_3_port);
   S4_4 : FA_X1 port map( A => ab_7_4_port, B => CARRYB_6_4_port, CI => 
                           SUMB_6_5_port, CO => CARRYB_7_4_port, S => 
                           SUMB_7_4_port);
   S4_5 : FA_X1 port map( A => ab_7_5_port, B => CARRYB_6_5_port, CI => 
                           SUMB_6_6_port, CO => CARRYB_7_5_port, S => 
                           SUMB_7_5_port);
   S5_6 : FA_X1 port map( A => ab_7_6_port, B => CARRYB_6_6_port, CI => 
                           ab_6_7_port, CO => CARRYB_7_6_port, S => 
                           SUMB_7_6_port);
   S1_6_0 : FA_X1 port map( A => ab_6_0_port, B => CARRYB_5_0_port, CI => 
                           SUMB_5_1_port, CO => CARRYB_6_0_port, S => A1_4_port
                           );
   S2_6_1 : FA_X1 port map( A => ab_6_1_port, B => CARRYB_5_1_port, CI => 
                           SUMB_5_2_port, CO => CARRYB_6_1_port, S => 
                           SUMB_6_1_port);
   S2_6_2 : FA_X1 port map( A => ab_6_2_port, B => CARRYB_5_2_port, CI => 
                           SUMB_5_3_port, CO => CARRYB_6_2_port, S => 
                           SUMB_6_2_port);
   S2_6_3 : FA_X1 port map( A => ab_6_3_port, B => CARRYB_5_3_port, CI => 
                           SUMB_5_4_port, CO => CARRYB_6_3_port, S => 
                           SUMB_6_3_port);
   S2_6_4 : FA_X1 port map( A => ab_6_4_port, B => CARRYB_5_4_port, CI => 
                           SUMB_5_5_port, CO => CARRYB_6_4_port, S => 
                           SUMB_6_4_port);
   S2_6_5 : FA_X1 port map( A => ab_6_5_port, B => CARRYB_5_5_port, CI => 
                           SUMB_5_6_port, CO => CARRYB_6_5_port, S => 
                           SUMB_6_5_port);
   S3_6_6 : FA_X1 port map( A => ab_6_6_port, B => CARRYB_5_6_port, CI => 
                           ab_5_7_port, CO => CARRYB_6_6_port, S => 
                           SUMB_6_6_port);
   S1_5_0 : FA_X1 port map( A => ab_5_0_port, B => CARRYB_4_0_port, CI => 
                           SUMB_4_1_port, CO => CARRYB_5_0_port, S => A1_3_port
                           );
   S2_5_1 : FA_X1 port map( A => ab_5_1_port, B => CARRYB_4_1_port, CI => 
                           SUMB_4_2_port, CO => CARRYB_5_1_port, S => 
                           SUMB_5_1_port);
   S2_5_2 : FA_X1 port map( A => ab_5_2_port, B => CARRYB_4_2_port, CI => 
                           SUMB_4_3_port, CO => CARRYB_5_2_port, S => 
                           SUMB_5_2_port);
   S2_5_3 : FA_X1 port map( A => ab_5_3_port, B => CARRYB_4_3_port, CI => 
                           SUMB_4_4_port, CO => CARRYB_5_3_port, S => 
                           SUMB_5_3_port);
   S2_5_4 : FA_X1 port map( A => ab_5_4_port, B => CARRYB_4_4_port, CI => 
                           SUMB_4_5_port, CO => CARRYB_5_4_port, S => 
                           SUMB_5_4_port);
   S2_5_5 : FA_X1 port map( A => ab_5_5_port, B => CARRYB_4_5_port, CI => 
                           SUMB_4_6_port, CO => CARRYB_5_5_port, S => 
                           SUMB_5_5_port);
   S3_5_6 : FA_X1 port map( A => ab_5_6_port, B => CARRYB_4_6_port, CI => 
                           ab_4_7_port, CO => CARRYB_5_6_port, S => 
                           SUMB_5_6_port);
   S1_4_0 : FA_X1 port map( A => ab_4_0_port, B => CARRYB_3_0_port, CI => 
                           SUMB_3_1_port, CO => CARRYB_4_0_port, S => A1_2_port
                           );
   S2_4_1 : FA_X1 port map( A => ab_4_1_port, B => CARRYB_3_1_port, CI => 
                           SUMB_3_2_port, CO => CARRYB_4_1_port, S => 
                           SUMB_4_1_port);
   S2_4_2 : FA_X1 port map( A => ab_4_2_port, B => CARRYB_3_2_port, CI => 
                           SUMB_3_3_port, CO => CARRYB_4_2_port, S => 
                           SUMB_4_2_port);
   S2_4_3 : FA_X1 port map( A => ab_4_3_port, B => CARRYB_3_3_port, CI => 
                           SUMB_3_4_port, CO => CARRYB_4_3_port, S => 
                           SUMB_4_3_port);
   S2_4_4 : FA_X1 port map( A => ab_4_4_port, B => CARRYB_3_4_port, CI => 
                           SUMB_3_5_port, CO => CARRYB_4_4_port, S => 
                           SUMB_4_4_port);
   S2_4_5 : FA_X1 port map( A => ab_4_5_port, B => CARRYB_3_5_port, CI => 
                           SUMB_3_6_port, CO => CARRYB_4_5_port, S => 
                           SUMB_4_5_port);
   S3_4_6 : FA_X1 port map( A => ab_4_6_port, B => CARRYB_3_6_port, CI => 
                           ab_3_7_port, CO => CARRYB_4_6_port, S => 
                           SUMB_4_6_port);
   S1_3_0 : FA_X1 port map( A => ab_3_0_port, B => CARRYB_2_0_port, CI => 
                           SUMB_2_1_port, CO => CARRYB_3_0_port, S => A1_1_port
                           );
   S2_3_1 : FA_X1 port map( A => ab_3_1_port, B => CARRYB_2_1_port, CI => 
                           SUMB_2_2_port, CO => CARRYB_3_1_port, S => 
                           SUMB_3_1_port);
   S2_3_2 : FA_X1 port map( A => ab_3_2_port, B => CARRYB_2_2_port, CI => 
                           SUMB_2_3_port, CO => CARRYB_3_2_port, S => 
                           SUMB_3_2_port);
   S2_3_3 : FA_X1 port map( A => ab_3_3_port, B => CARRYB_2_3_port, CI => 
                           SUMB_2_4_port, CO => CARRYB_3_3_port, S => 
                           SUMB_3_3_port);
   S2_3_4 : FA_X1 port map( A => ab_3_4_port, B => CARRYB_2_4_port, CI => 
                           SUMB_2_5_port, CO => CARRYB_3_4_port, S => 
                           SUMB_3_4_port);
   S2_3_5 : FA_X1 port map( A => ab_3_5_port, B => CARRYB_2_5_port, CI => 
                           SUMB_2_6_port, CO => CARRYB_3_5_port, S => 
                           SUMB_3_5_port);
   S3_3_6 : FA_X1 port map( A => ab_3_6_port, B => CARRYB_2_6_port, CI => 
                           ab_2_7_port, CO => CARRYB_3_6_port, S => 
                           SUMB_3_6_port);
   S1_2_0 : FA_X1 port map( A => ab_2_0_port, B => n7, CI => n14, CO => 
                           CARRYB_2_0_port, S => A1_0_port);
   S2_2_1 : FA_X1 port map( A => ab_2_1_port, B => n6, CI => n13, CO => 
                           CARRYB_2_1_port, S => SUMB_2_1_port);
   S2_2_2 : FA_X1 port map( A => ab_2_2_port, B => n5, CI => n12, CO => 
                           CARRYB_2_2_port, S => SUMB_2_2_port);
   S2_2_3 : FA_X1 port map( A => ab_2_3_port, B => n4, CI => n11, CO => 
                           CARRYB_2_3_port, S => SUMB_2_3_port);
   S2_2_4 : FA_X1 port map( A => ab_2_4_port, B => n3, CI => n10, CO => 
                           CARRYB_2_4_port, S => SUMB_2_4_port);
   S2_2_5 : FA_X1 port map( A => ab_2_5_port, B => n2, CI => n9, CO => 
                           CARRYB_2_5_port, S => SUMB_2_5_port);
   S3_2_6 : FA_X1 port map( A => ab_2_6_port, B => n8, CI => ab_1_7_port, CO =>
                           CARRYB_2_6_port, S => SUMB_2_6_port);
   FS_1 : shift_pow2_N8_1_DW01_add_0 port map( A(13) => n46, A(12) => n17, 
                           A(11) => n21, A(10) => n19, A(9) => n22, A(8) => n27
                           , A(7) => n20, A(6) => n18, A(5) => SUMB_7_0_port, 
                           A(4) => A1_4_port, A(3) => A1_3_port, A(2) => 
                           A1_2_port, A(1) => A1_1_port, A(0) => A1_0_port, 
                           B(13) => n15, B(12) => n28, B(11) => n25, B(10) => 
                           n23, B(9) => n26, B(8) => n29, B(7) => n24, B(6) => 
                           n46, B(5) => n47, B(4) => n47, B(3) => n47, B(2) => 
                           n47, B(1) => n47, B(0) => X_Logic0_port, CI => 
                           X_Logic0_port, SUM(13) => PRODUCT(15), SUM(12) => 
                           PRODUCT(14), SUM(11) => PRODUCT(13), SUM(10) => 
                           PRODUCT(12), SUM(9) => PRODUCT(11), SUM(8) => 
                           PRODUCT(10), SUM(7) => PRODUCT(9), SUM(6) => 
                           PRODUCT(8), SUM(5) => PRODUCT(7), SUM(4) => 
                           PRODUCT(6), SUM(3) => PRODUCT(5), SUM(2) => 
                           PRODUCT(4), SUM(1) => PRODUCT(3), SUM(0) => 
                           PRODUCT(2), CO => n_1095);
   U2 : INV_X1 port map( A => B(4), ZN => n35);
   U3 : INV_X1 port map( A => B(5), ZN => n34);
   U4 : INV_X1 port map( A => B(6), ZN => n33);
   U5 : INV_X1 port map( A => B(7), ZN => n30);
   U6 : AND2_X1 port map( A1 => ab_0_6_port, A2 => ab_1_5_port, ZN => n2);
   U7 : AND2_X1 port map( A1 => ab_0_5_port, A2 => ab_1_4_port, ZN => n3);
   U8 : AND2_X1 port map( A1 => ab_0_4_port, A2 => ab_1_3_port, ZN => n4);
   U9 : AND2_X1 port map( A1 => ab_0_3_port, A2 => ab_1_2_port, ZN => n5);
   U10 : AND2_X1 port map( A1 => ab_0_2_port, A2 => ab_1_1_port, ZN => n6);
   U11 : AND2_X1 port map( A1 => ab_0_1_port, A2 => ab_1_0_port, ZN => n7);
   U12 : AND2_X1 port map( A1 => ab_0_7_port, A2 => ab_1_6_port, ZN => n8);
   U13 : XOR2_X1 port map( A => ab_1_6_port, B => ab_0_7_port, Z => n9);
   U14 : XOR2_X1 port map( A => ab_1_5_port, B => ab_0_6_port, Z => n10);
   U15 : XOR2_X1 port map( A => ab_1_4_port, B => ab_0_5_port, Z => n11);
   U16 : XOR2_X1 port map( A => ab_1_3_port, B => ab_0_4_port, Z => n12);
   U17 : XOR2_X1 port map( A => ab_1_2_port, B => ab_0_3_port, Z => n13);
   U18 : XOR2_X1 port map( A => ab_1_1_port, B => ab_0_2_port, Z => n14);
   U19 : AND2_X1 port map( A1 => CARRYB_7_6_port, A2 => ab_7_7_port, ZN => n15)
                           ;
   U20 : XOR2_X1 port map( A => ab_1_0_port, B => ab_0_1_port, Z => PRODUCT(1))
                           ;
   U21 : XOR2_X1 port map( A => CARRYB_7_6_port, B => ab_7_7_port, Z => n17);
   U22 : XOR2_X1 port map( A => CARRYB_7_0_port, B => SUMB_7_1_port, Z => n18);
   U23 : XOR2_X1 port map( A => CARRYB_7_4_port, B => SUMB_7_5_port, Z => n19);
   U24 : XOR2_X1 port map( A => CARRYB_7_1_port, B => SUMB_7_2_port, Z => n20);
   U25 : XOR2_X1 port map( A => CARRYB_7_5_port, B => SUMB_7_6_port, Z => n21);
   U26 : XOR2_X1 port map( A => CARRYB_7_3_port, B => SUMB_7_4_port, Z => n22);
   U27 : AND2_X1 port map( A1 => CARRYB_7_3_port, A2 => SUMB_7_4_port, ZN => 
                           n23);
   U28 : AND2_X1 port map( A1 => CARRYB_7_0_port, A2 => SUMB_7_1_port, ZN => 
                           n24);
   U29 : AND2_X1 port map( A1 => CARRYB_7_4_port, A2 => SUMB_7_5_port, ZN => 
                           n25);
   U30 : AND2_X1 port map( A1 => CARRYB_7_2_port, A2 => SUMB_7_3_port, ZN => 
                           n26);
   U31 : XOR2_X1 port map( A => CARRYB_7_2_port, B => SUMB_7_3_port, Z => n27);
   U32 : AND2_X1 port map( A1 => CARRYB_7_5_port, A2 => SUMB_7_6_port, ZN => 
                           n28);
   U33 : AND2_X1 port map( A1 => CARRYB_7_1_port, A2 => SUMB_7_2_port, ZN => 
                           n29);
   U34 : INV_X1 port map( A => B(2), ZN => n32);
   U35 : INV_X1 port map( A => B(1), ZN => n36);
   U36 : INV_X1 port map( A => B(3), ZN => n31);
   U37 : INV_X1 port map( A => B(0), ZN => n37);
   U38 : INV_X1 port map( A => A(7), ZN => n38);
   U39 : INV_X1 port map( A => A(0), ZN => n45);
   U40 : INV_X1 port map( A => A(1), ZN => n44);
   U41 : INV_X1 port map( A => A(2), ZN => n43);
   U42 : INV_X1 port map( A => A(3), ZN => n42);
   U43 : INV_X1 port map( A => A(4), ZN => n41);
   U44 : INV_X1 port map( A => A(5), ZN => n40);
   U45 : INV_X1 port map( A => A(6), ZN => n39);
   n46 <= '0';
   U47 : NOR2_X1 port map( A1 => n38, A2 => n30, ZN => ab_7_7_port);
   U48 : NOR2_X1 port map( A1 => n38, A2 => n33, ZN => ab_7_6_port);
   U49 : NOR2_X1 port map( A1 => n38, A2 => n34, ZN => ab_7_5_port);
   U50 : NOR2_X1 port map( A1 => n38, A2 => n35, ZN => ab_7_4_port);
   U51 : NOR2_X1 port map( A1 => n38, A2 => n31, ZN => ab_7_3_port);
   U52 : NOR2_X1 port map( A1 => n38, A2 => n32, ZN => ab_7_2_port);
   U53 : NOR2_X1 port map( A1 => n38, A2 => n36, ZN => ab_7_1_port);
   U54 : NOR2_X1 port map( A1 => n38, A2 => n37, ZN => ab_7_0_port);
   U55 : NOR2_X1 port map( A1 => n30, A2 => n39, ZN => ab_6_7_port);
   U56 : NOR2_X1 port map( A1 => n33, A2 => n39, ZN => ab_6_6_port);
   U57 : NOR2_X1 port map( A1 => n34, A2 => n39, ZN => ab_6_5_port);
   U58 : NOR2_X1 port map( A1 => n35, A2 => n39, ZN => ab_6_4_port);
   U59 : NOR2_X1 port map( A1 => n31, A2 => n39, ZN => ab_6_3_port);
   U60 : NOR2_X1 port map( A1 => n32, A2 => n39, ZN => ab_6_2_port);
   U61 : NOR2_X1 port map( A1 => n36, A2 => n39, ZN => ab_6_1_port);
   U62 : NOR2_X1 port map( A1 => n37, A2 => n39, ZN => ab_6_0_port);
   U63 : NOR2_X1 port map( A1 => n30, A2 => n40, ZN => ab_5_7_port);
   U64 : NOR2_X1 port map( A1 => n33, A2 => n40, ZN => ab_5_6_port);
   U65 : NOR2_X1 port map( A1 => n34, A2 => n40, ZN => ab_5_5_port);
   U66 : NOR2_X1 port map( A1 => n35, A2 => n40, ZN => ab_5_4_port);
   U67 : NOR2_X1 port map( A1 => n31, A2 => n40, ZN => ab_5_3_port);
   U68 : NOR2_X1 port map( A1 => n32, A2 => n40, ZN => ab_5_2_port);
   U69 : NOR2_X1 port map( A1 => n36, A2 => n40, ZN => ab_5_1_port);
   U70 : NOR2_X1 port map( A1 => n37, A2 => n40, ZN => ab_5_0_port);
   U71 : NOR2_X1 port map( A1 => n30, A2 => n41, ZN => ab_4_7_port);
   U72 : NOR2_X1 port map( A1 => n33, A2 => n41, ZN => ab_4_6_port);
   U73 : NOR2_X1 port map( A1 => n34, A2 => n41, ZN => ab_4_5_port);
   U74 : NOR2_X1 port map( A1 => n35, A2 => n41, ZN => ab_4_4_port);
   U75 : NOR2_X1 port map( A1 => n31, A2 => n41, ZN => ab_4_3_port);
   U76 : NOR2_X1 port map( A1 => n32, A2 => n41, ZN => ab_4_2_port);
   U77 : NOR2_X1 port map( A1 => n36, A2 => n41, ZN => ab_4_1_port);
   U78 : NOR2_X1 port map( A1 => n37, A2 => n41, ZN => ab_4_0_port);
   U79 : NOR2_X1 port map( A1 => n30, A2 => n42, ZN => ab_3_7_port);
   U80 : NOR2_X1 port map( A1 => n33, A2 => n42, ZN => ab_3_6_port);
   U81 : NOR2_X1 port map( A1 => n34, A2 => n42, ZN => ab_3_5_port);
   U82 : NOR2_X1 port map( A1 => n35, A2 => n42, ZN => ab_3_4_port);
   U83 : NOR2_X1 port map( A1 => n31, A2 => n42, ZN => ab_3_3_port);
   U84 : NOR2_X1 port map( A1 => n32, A2 => n42, ZN => ab_3_2_port);
   U85 : NOR2_X1 port map( A1 => n36, A2 => n42, ZN => ab_3_1_port);
   U86 : NOR2_X1 port map( A1 => n37, A2 => n42, ZN => ab_3_0_port);
   U87 : NOR2_X1 port map( A1 => n30, A2 => n43, ZN => ab_2_7_port);
   U88 : NOR2_X1 port map( A1 => n33, A2 => n43, ZN => ab_2_6_port);
   U89 : NOR2_X1 port map( A1 => n34, A2 => n43, ZN => ab_2_5_port);
   U90 : NOR2_X1 port map( A1 => n35, A2 => n43, ZN => ab_2_4_port);
   U91 : NOR2_X1 port map( A1 => n31, A2 => n43, ZN => ab_2_3_port);
   U92 : NOR2_X1 port map( A1 => n32, A2 => n43, ZN => ab_2_2_port);
   U93 : NOR2_X1 port map( A1 => n36, A2 => n43, ZN => ab_2_1_port);
   U94 : NOR2_X1 port map( A1 => n37, A2 => n43, ZN => ab_2_0_port);
   U95 : NOR2_X1 port map( A1 => n30, A2 => n44, ZN => ab_1_7_port);
   U96 : NOR2_X1 port map( A1 => n33, A2 => n44, ZN => ab_1_6_port);
   U97 : NOR2_X1 port map( A1 => n34, A2 => n44, ZN => ab_1_5_port);
   U98 : NOR2_X1 port map( A1 => n35, A2 => n44, ZN => ab_1_4_port);
   U99 : NOR2_X1 port map( A1 => n31, A2 => n44, ZN => ab_1_3_port);
   U100 : NOR2_X1 port map( A1 => n32, A2 => n44, ZN => ab_1_2_port);
   U101 : NOR2_X1 port map( A1 => n36, A2 => n44, ZN => ab_1_1_port);
   U102 : NOR2_X1 port map( A1 => n37, A2 => n44, ZN => ab_1_0_port);
   U103 : NOR2_X1 port map( A1 => n30, A2 => n45, ZN => ab_0_7_port);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n45, ZN => ab_0_6_port);
   U105 : NOR2_X1 port map( A1 => n34, A2 => n45, ZN => ab_0_5_port);
   U106 : NOR2_X1 port map( A1 => n35, A2 => n45, ZN => ab_0_4_port);
   U107 : NOR2_X1 port map( A1 => n31, A2 => n45, ZN => ab_0_3_port);
   U108 : NOR2_X1 port map( A1 => n32, A2 => n45, ZN => ab_0_2_port);
   U109 : NOR2_X1 port map( A1 => n36, A2 => n45, ZN => ab_0_1_port);
   U110 : NOR2_X1 port map( A1 => n37, A2 => n45, ZN => PRODUCT(0));
   n47 <= '0';

end SYN_csa;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_0_DW01_inc_0_DW01_inc_7 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end complementor_N16_0_DW01_inc_0_DW01_inc_7;

architecture SYN_rpl of complementor_N16_0_DW01_inc_0_DW01_inc_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port : 
      std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_7_DW01_inc_0_DW01_inc_6 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end complementor_N16_7_DW01_inc_0_DW01_inc_6;

architecture SYN_rpl of complementor_N16_7_DW01_inc_0_DW01_inc_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port : 
      std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_6_DW01_inc_0_DW01_inc_5 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end complementor_N16_6_DW01_inc_0_DW01_inc_5;

architecture SYN_rpl of complementor_N16_6_DW01_inc_0_DW01_inc_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port : 
      std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_5_DW01_inc_0_DW01_inc_4 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end complementor_N16_5_DW01_inc_0_DW01_inc_4;

architecture SYN_rpl of complementor_N16_5_DW01_inc_0_DW01_inc_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port : 
      std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_4_DW01_inc_0_DW01_inc_3 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end complementor_N16_4_DW01_inc_0_DW01_inc_3;

architecture SYN_rpl of complementor_N16_4_DW01_inc_0_DW01_inc_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port : 
      std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_3_DW01_inc_0_DW01_inc_2 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end complementor_N16_3_DW01_inc_0_DW01_inc_2;

architecture SYN_rpl of complementor_N16_3_DW01_inc_0_DW01_inc_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port : 
      std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_2_DW01_inc_0_DW01_inc_1 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end complementor_N16_2_DW01_inc_0_DW01_inc_1;

architecture SYN_rpl of complementor_N16_2_DW01_inc_0_DW01_inc_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port : 
      std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_1_DW01_inc_0 is

   port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector (15
         downto 0));

end complementor_N16_1_DW01_inc_0;

architecture SYN_rpl of complementor_N16_1_DW01_inc_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port : 
      std_logic;

begin
   
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_15_port, B => A(15), Z => SUM(15));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2015 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2015;

architecture SYN_ARCHBEH of FA_2015 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2014 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2014;

architecture SYN_ARCHBEH of FA_2014 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2013 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2013;

architecture SYN_ARCHBEH of FA_2013 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2012 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2012;

architecture SYN_ARCHBEH of FA_2012 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2011 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2011;

architecture SYN_ARCHBEH of FA_2011 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2010 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2010;

architecture SYN_ARCHBEH of FA_2010 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2009 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2009;

architecture SYN_ARCHBEH of FA_2009 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2008 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2008;

architecture SYN_ARCHBEH of FA_2008 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2007 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2007;

architecture SYN_ARCHBEH of FA_2007 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2006 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2006;

architecture SYN_ARCHBEH of FA_2006 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2005 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2005;

architecture SYN_ARCHBEH of FA_2005 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2004 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2004;

architecture SYN_ARCHBEH of FA_2004 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2003 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2003;

architecture SYN_ARCHBEH of FA_2003 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2002 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2002;

architecture SYN_ARCHBEH of FA_2002 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2001 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2001;

architecture SYN_ARCHBEH of FA_2001 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_2000 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2000;

architecture SYN_ARCHBEH of FA_2000 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1999 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1999;

architecture SYN_ARCHBEH of FA_1999 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1998 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1998;

architecture SYN_ARCHBEH of FA_1998 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1997 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1997;

architecture SYN_ARCHBEH of FA_1997 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1996 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1996;

architecture SYN_ARCHBEH of FA_1996 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1995 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1995;

architecture SYN_ARCHBEH of FA_1995 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1994 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1994;

architecture SYN_ARCHBEH of FA_1994 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1993 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1993;

architecture SYN_ARCHBEH of FA_1993 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1992 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1992;

architecture SYN_ARCHBEH of FA_1992 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1991 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1991;

architecture SYN_ARCHBEH of FA_1991 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1990 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1990;

architecture SYN_ARCHBEH of FA_1990 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1989 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1989;

architecture SYN_ARCHBEH of FA_1989 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1988 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1988;

architecture SYN_ARCHBEH of FA_1988 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1987 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1987;

architecture SYN_ARCHBEH of FA_1987 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1986 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1986;

architecture SYN_ARCHBEH of FA_1986 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1985 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1985;

architecture SYN_ARCHBEH of FA_1985 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1984 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1984;

architecture SYN_ARCHBEH of FA_1984 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1983 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1983;

architecture SYN_ARCHBEH of FA_1983 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1982 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1982;

architecture SYN_ARCHBEH of FA_1982 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1981 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1981;

architecture SYN_ARCHBEH of FA_1981 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1980 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1980;

architecture SYN_ARCHBEH of FA_1980 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1979 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1979;

architecture SYN_ARCHBEH of FA_1979 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1978 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1978;

architecture SYN_ARCHBEH of FA_1978 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1977 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1977;

architecture SYN_ARCHBEH of FA_1977 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1976 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1976;

architecture SYN_ARCHBEH of FA_1976 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1975 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1975;

architecture SYN_ARCHBEH of FA_1975 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1974 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1974;

architecture SYN_ARCHBEH of FA_1974 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1973 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1973;

architecture SYN_ARCHBEH of FA_1973 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1972 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1972;

architecture SYN_ARCHBEH of FA_1972 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1971 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1971;

architecture SYN_ARCHBEH of FA_1971 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1970 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1970;

architecture SYN_ARCHBEH of FA_1970 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1969 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1969;

architecture SYN_ARCHBEH of FA_1969 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1968 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1968;

architecture SYN_ARCHBEH of FA_1968 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1967 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1967;

architecture SYN_ARCHBEH of FA_1967 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1966 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1966;

architecture SYN_ARCHBEH of FA_1966 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1965 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1965;

architecture SYN_ARCHBEH of FA_1965 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1964 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1964;

architecture SYN_ARCHBEH of FA_1964 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1963 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1963;

architecture SYN_ARCHBEH of FA_1963 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1962 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1962;

architecture SYN_ARCHBEH of FA_1962 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1961 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1961;

architecture SYN_ARCHBEH of FA_1961 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1960 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1960;

architecture SYN_ARCHBEH of FA_1960 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1959 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1959;

architecture SYN_ARCHBEH of FA_1959 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1958 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1958;

architecture SYN_ARCHBEH of FA_1958 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1957 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1957;

architecture SYN_ARCHBEH of FA_1957 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1956 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1956;

architecture SYN_ARCHBEH of FA_1956 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1955 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1955;

architecture SYN_ARCHBEH of FA_1955 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1954 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1954;

architecture SYN_ARCHBEH of FA_1954 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1953 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1953;

architecture SYN_ARCHBEH of FA_1953 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1952 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1952;

architecture SYN_ARCHBEH of FA_1952 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1951 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1951;

architecture SYN_ARCHBEH of FA_1951 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1950 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1950;

architecture SYN_ARCHBEH of FA_1950 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1949 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1949;

architecture SYN_ARCHBEH of FA_1949 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1948 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1948;

architecture SYN_ARCHBEH of FA_1948 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1947 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1947;

architecture SYN_ARCHBEH of FA_1947 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1946 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1946;

architecture SYN_ARCHBEH of FA_1946 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1945 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1945;

architecture SYN_ARCHBEH of FA_1945 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1944 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1944;

architecture SYN_ARCHBEH of FA_1944 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1943 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1943;

architecture SYN_ARCHBEH of FA_1943 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1942 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1942;

architecture SYN_ARCHBEH of FA_1942 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1941 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1941;

architecture SYN_ARCHBEH of FA_1941 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1940 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1940;

architecture SYN_ARCHBEH of FA_1940 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1939 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1939;

architecture SYN_ARCHBEH of FA_1939 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1938 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1938;

architecture SYN_ARCHBEH of FA_1938 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1937 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1937;

architecture SYN_ARCHBEH of FA_1937 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1936 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1936;

architecture SYN_ARCHBEH of FA_1936 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1935 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1935;

architecture SYN_ARCHBEH of FA_1935 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1934 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1934;

architecture SYN_ARCHBEH of FA_1934 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1933 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1933;

architecture SYN_ARCHBEH of FA_1933 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1932 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1932;

architecture SYN_ARCHBEH of FA_1932 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1931 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1931;

architecture SYN_ARCHBEH of FA_1931 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1930 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1930;

architecture SYN_ARCHBEH of FA_1930 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1929 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1929;

architecture SYN_ARCHBEH of FA_1929 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1928 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1928;

architecture SYN_ARCHBEH of FA_1928 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1927 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1927;

architecture SYN_ARCHBEH of FA_1927 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1926 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1926;

architecture SYN_ARCHBEH of FA_1926 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1925 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1925;

architecture SYN_ARCHBEH of FA_1925 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1924 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1924;

architecture SYN_ARCHBEH of FA_1924 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1923 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1923;

architecture SYN_ARCHBEH of FA_1923 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1922 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1922;

architecture SYN_ARCHBEH of FA_1922 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1921 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1921;

architecture SYN_ARCHBEH of FA_1921 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_251 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_251;

architecture SYN_ARCHSTRUCT of muxN1_N4_251 is

   component mux21_8169
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8170
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8171
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8172
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8172 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8171 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8170 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8169 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_250 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_250;

architecture SYN_ARCHSTRUCT of muxN1_N4_250 is

   component mux21_8165
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8166
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8167
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8168
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8168 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8167 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8166 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8165 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_249 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_249;

architecture SYN_ARCHSTRUCT of muxN1_N4_249 is

   component mux21_8161
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8162
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8163
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8164
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8164 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8163 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8162 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8161 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_248 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_248;

architecture SYN_ARCHSTRUCT of muxN1_N4_248 is

   component mux21_8157
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8158
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8159
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8160
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8160 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8159 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8158 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8157 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_247 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_247;

architecture SYN_ARCHSTRUCT of muxN1_N4_247 is

   component mux21_8153
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8154
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8155
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8156
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8156 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8155 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8154 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8153 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_246 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_246;

architecture SYN_ARCHSTRUCT of muxN1_N4_246 is

   component mux21_8149
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8150
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8151
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8152
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8152 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8151 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8150 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8149 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_245 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_245;

architecture SYN_ARCHSTRUCT of muxN1_N4_245 is

   component mux21_8145
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8146
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8147
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8148
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8148 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8147 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8146 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8145 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_244 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_244;

architecture SYN_ARCHSTRUCT of muxN1_N4_244 is

   component mux21_8141
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8142
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8143
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8144
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8144 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8143 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8142 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8141 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_243 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_243;

architecture SYN_ARCHSTRUCT of muxN1_N4_243 is

   component mux21_8137
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8138
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8139
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8140
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8140 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8139 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8138 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8137 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_242 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_242;

architecture SYN_ARCHSTRUCT of muxN1_N4_242 is

   component mux21_8133
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8134
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8135
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8136
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8136 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8135 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8134 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8133 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_241 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_241;

architecture SYN_ARCHSTRUCT of muxN1_N4_241 is

   component mux21_8129
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8130
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8131
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8132
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8132 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8131 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8130 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8129 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_503 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_503;

architecture SYN_ARCHSTRUCT of RCA_N4_503 is

   component FA_2009
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2010
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2011
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2012
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_2012 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_2011 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_2010 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_2009 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_502 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_502;

architecture SYN_ARCHSTRUCT of RCA_N4_502 is

   component FA_2005
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2006
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2007
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2008
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_2008 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_2007 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_2006 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_2005 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_501 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_501;

architecture SYN_ARCHSTRUCT of RCA_N4_501 is

   component FA_2001
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2002
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2003
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2004
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_2004 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_2003 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_2002 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_2001 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_500 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_500;

architecture SYN_ARCHSTRUCT of RCA_N4_500 is

   component FA_1997
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1998
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1999
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2000
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_2000 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1999 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1998 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1997 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_499 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_499;

architecture SYN_ARCHSTRUCT of RCA_N4_499 is

   component FA_1993
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1994
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1995
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1996
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1996 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1995 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1994 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1993 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_498 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_498;

architecture SYN_ARCHSTRUCT of RCA_N4_498 is

   component FA_1989
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1990
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1991
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1992
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1992 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1991 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1990 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1989 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_497 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_497;

architecture SYN_ARCHSTRUCT of RCA_N4_497 is

   component FA_1985
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1986
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1987
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1988
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1988 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1987 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1986 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1985 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_496 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_496;

architecture SYN_ARCHSTRUCT of RCA_N4_496 is

   component FA_1981
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1982
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1983
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1984
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1984 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1983 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1982 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1981 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_495 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_495;

architecture SYN_ARCHSTRUCT of RCA_N4_495 is

   component FA_1977
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1978
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1979
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1980
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1980 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1979 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1978 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1977 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_494 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_494;

architecture SYN_ARCHSTRUCT of RCA_N4_494 is

   component FA_1973
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1974
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1975
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1976
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1976 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1975 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1974 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1973 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_493 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_493;

architecture SYN_ARCHSTRUCT of RCA_N4_493 is

   component FA_1969
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1970
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1971
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1972
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1972 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1971 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1970 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1969 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_492 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_492;

architecture SYN_ARCHSTRUCT of RCA_N4_492 is

   component FA_1965
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1966
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1967
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1968
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1968 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1967 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1966 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1965 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_491 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_491;

architecture SYN_ARCHSTRUCT of RCA_N4_491 is

   component FA_1961
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1962
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1963
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1964
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1964 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1963 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1962 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1961 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_490 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_490;

architecture SYN_ARCHSTRUCT of RCA_N4_490 is

   component FA_1957
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1958
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1959
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1960
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1960 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1959 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1958 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1957 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_489 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_489;

architecture SYN_ARCHSTRUCT of RCA_N4_489 is

   component FA_1953
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1954
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1955
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1956
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1956 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1955 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1954 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1953 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_488 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_488;

architecture SYN_ARCHSTRUCT of RCA_N4_488 is

   component FA_1949
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1950
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1951
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1952
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1952 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1951 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1950 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1949 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_487 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_487;

architecture SYN_ARCHSTRUCT of RCA_N4_487 is

   component FA_1945
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1946
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1947
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1948
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1948 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1947 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1946 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1945 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_486 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_486;

architecture SYN_ARCHSTRUCT of RCA_N4_486 is

   component FA_1941
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1942
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1943
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1944
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1944 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1943 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1942 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1941 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_485 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_485;

architecture SYN_ARCHSTRUCT of RCA_N4_485 is

   component FA_1937
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1938
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1939
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1940
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1940 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1939 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1938 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1937 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_484 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_484;

architecture SYN_ARCHSTRUCT of RCA_N4_484 is

   component FA_1933
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1934
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1935
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1936
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1936 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1935 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1934 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1933 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_483 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_483;

architecture SYN_ARCHSTRUCT of RCA_N4_483 is

   component FA_1929
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1930
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1931
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1932
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1932 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1931 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1930 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1929 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_482 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_482;

architecture SYN_ARCHSTRUCT of RCA_N4_482 is

   component FA_1925
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1926
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1927
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1928
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1928 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1927 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1926 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1925 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_481 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_481;

architecture SYN_ARCHSTRUCT of RCA_N4_481 is

   component FA_1921
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1922
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1923
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1924
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1924 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1923 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1922 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1921 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_977 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_977;

architecture SYN_ARCHDATAFLOW of pg_block_977 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_976 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_976;

architecture SYN_ARCHDATAFLOW of pg_block_976 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_975 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_975;

architecture SYN_ARCHDATAFLOW of pg_block_975 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_974 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_974;

architecture SYN_ARCHDATAFLOW of pg_block_974 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_973 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_973;

architecture SYN_ARCHDATAFLOW of pg_block_973 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_972 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_972;

architecture SYN_ARCHDATAFLOW of pg_block_972 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_971 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_971;

architecture SYN_ARCHDATAFLOW of pg_block_971 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_970 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_970;

architecture SYN_ARCHDATAFLOW of pg_block_970 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_969 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_969;

architecture SYN_ARCHDATAFLOW of pg_block_969 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_968 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_968;

architecture SYN_ARCHDATAFLOW of pg_block_968 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_967 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_967;

architecture SYN_ARCHDATAFLOW of pg_block_967 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_966 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_966;

architecture SYN_ARCHDATAFLOW of pg_block_966 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_965 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_965;

architecture SYN_ARCHDATAFLOW of pg_block_965 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_964 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_964;

architecture SYN_ARCHDATAFLOW of pg_block_964 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_963 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_963;

architecture SYN_ARCHDATAFLOW of pg_block_963 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_962 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_962;

architecture SYN_ARCHDATAFLOW of pg_block_962 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_961 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_961;

architecture SYN_ARCHDATAFLOW of pg_block_961 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_960 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_960;

architecture SYN_ARCHDATAFLOW of pg_block_960 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_959 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_959;

architecture SYN_ARCHDATAFLOW of pg_block_959 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_958 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_958;

architecture SYN_ARCHDATAFLOW of pg_block_958 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_957 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_957;

architecture SYN_ARCHDATAFLOW of pg_block_957 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_956 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_956;

architecture SYN_ARCHDATAFLOW of pg_block_956 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_955 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_955;

architecture SYN_ARCHDATAFLOW of pg_block_955 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_954 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_954;

architecture SYN_ARCHDATAFLOW of pg_block_954 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_953 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_953;

architecture SYN_ARCHDATAFLOW of pg_block_953 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_952 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_952;

architecture SYN_ARCHDATAFLOW of pg_block_952 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_951 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_951;

architecture SYN_ARCHDATAFLOW of pg_block_951 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_950 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_950;

architecture SYN_ARCHDATAFLOW of pg_block_950 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_949 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_949;

architecture SYN_ARCHDATAFLOW of pg_block_949 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_948 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_948;

architecture SYN_ARCHDATAFLOW of pg_block_948 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_947 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_947;

architecture SYN_ARCHDATAFLOW of pg_block_947 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_946 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_946;

architecture SYN_ARCHDATAFLOW of pg_block_946 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_269 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_269;

architecture SYN_ARCHDATAFLOW of g_block_269 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_268 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_268;

architecture SYN_ARCHDATAFLOW of g_block_268 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_267 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_267;

architecture SYN_ARCHDATAFLOW of g_block_267 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_266 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_266;

architecture SYN_ARCHDATAFLOW of g_block_266 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_265 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_265;

architecture SYN_ARCHDATAFLOW of g_block_265 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_264 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_264;

architecture SYN_ARCHDATAFLOW of g_block_264 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_263 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_263;

architecture SYN_ARCHDATAFLOW of g_block_263 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_262 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_262;

architecture SYN_ARCHDATAFLOW of g_block_262 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_261 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_261;

architecture SYN_ARCHDATAFLOW of g_block_261 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_260 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_260;

architecture SYN_ARCHDATAFLOW of g_block_260 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_259 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_259;

architecture SYN_ARCHDATAFLOW of g_block_259 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_258 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_258;

architecture SYN_ARCHDATAFLOW of g_block_258 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_257 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_257;

architecture SYN_ARCHDATAFLOW of g_block_257 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_256 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_256;

architecture SYN_ARCHDATAFLOW of g_block_256 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25871 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25871;

architecture SYN_ARCHBEH of nd2_25871 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25870 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25870;

architecture SYN_ARCHBEH of nd2_25870 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25869 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25869;

architecture SYN_ARCHBEH of nd2_25869 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25868 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25868;

architecture SYN_ARCHBEH of nd2_25868 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25867 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25867;

architecture SYN_ARCHBEH of nd2_25867 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25866 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25866;

architecture SYN_ARCHBEH of nd2_25866 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25865 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25865;

architecture SYN_ARCHBEH of nd2_25865 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25864 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25864;

architecture SYN_ARCHBEH of nd2_25864 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25863 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25863;

architecture SYN_ARCHBEH of nd2_25863 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25862 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25862;

architecture SYN_ARCHBEH of nd2_25862 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25861 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25861;

architecture SYN_ARCHBEH of nd2_25861 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25860 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25860;

architecture SYN_ARCHBEH of nd2_25860 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25859 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25859;

architecture SYN_ARCHBEH of nd2_25859 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25858 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25858;

architecture SYN_ARCHBEH of nd2_25858 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25857 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25857;

architecture SYN_ARCHBEH of nd2_25857 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25856 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25856;

architecture SYN_ARCHBEH of nd2_25856 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25855 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25855;

architecture SYN_ARCHBEH of nd2_25855 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25854 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25854;

architecture SYN_ARCHBEH of nd2_25854 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25853 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25853;

architecture SYN_ARCHBEH of nd2_25853 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25852 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25852;

architecture SYN_ARCHBEH of nd2_25852 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25851 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25851;

architecture SYN_ARCHBEH of nd2_25851 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25850 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25850;

architecture SYN_ARCHBEH of nd2_25850 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25849 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25849;

architecture SYN_ARCHBEH of nd2_25849 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25848 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25848;

architecture SYN_ARCHBEH of nd2_25848 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25847 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25847;

architecture SYN_ARCHBEH of nd2_25847 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25846 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25846;

architecture SYN_ARCHBEH of nd2_25846 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25845 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25845;

architecture SYN_ARCHBEH of nd2_25845 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25844 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25844;

architecture SYN_ARCHBEH of nd2_25844 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25843 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25843;

architecture SYN_ARCHBEH of nd2_25843 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25842 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25842;

architecture SYN_ARCHBEH of nd2_25842 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25841 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25841;

architecture SYN_ARCHBEH of nd2_25841 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25840 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25840;

architecture SYN_ARCHBEH of nd2_25840 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25839 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25839;

architecture SYN_ARCHBEH of nd2_25839 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25838 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25838;

architecture SYN_ARCHBEH of nd2_25838 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25837 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25837;

architecture SYN_ARCHBEH of nd2_25837 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25836 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25836;

architecture SYN_ARCHBEH of nd2_25836 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25835 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25835;

architecture SYN_ARCHBEH of nd2_25835 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25834 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25834;

architecture SYN_ARCHBEH of nd2_25834 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25833 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25833;

architecture SYN_ARCHBEH of nd2_25833 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25832 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25832;

architecture SYN_ARCHBEH of nd2_25832 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25831 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25831;

architecture SYN_ARCHBEH of nd2_25831 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25830 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25830;

architecture SYN_ARCHBEH of nd2_25830 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25829 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25829;

architecture SYN_ARCHBEH of nd2_25829 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25828 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25828;

architecture SYN_ARCHBEH of nd2_25828 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25827 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25827;

architecture SYN_ARCHBEH of nd2_25827 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25826 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25826;

architecture SYN_ARCHBEH of nd2_25826 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25825 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25825;

architecture SYN_ARCHBEH of nd2_25825 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25824 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25824;

architecture SYN_ARCHBEH of nd2_25824 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25823 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25823;

architecture SYN_ARCHBEH of nd2_25823 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25822 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25822;

architecture SYN_ARCHBEH of nd2_25822 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25821 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25821;

architecture SYN_ARCHBEH of nd2_25821 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25820 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25820;

architecture SYN_ARCHBEH of nd2_25820 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25819 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25819;

architecture SYN_ARCHBEH of nd2_25819 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25818 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25818;

architecture SYN_ARCHBEH of nd2_25818 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25817 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25817;

architecture SYN_ARCHBEH of nd2_25817 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25816 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25816;

architecture SYN_ARCHBEH of nd2_25816 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25815 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25815;

architecture SYN_ARCHBEH of nd2_25815 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25814 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25814;

architecture SYN_ARCHBEH of nd2_25814 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25813 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25813;

architecture SYN_ARCHBEH of nd2_25813 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25812 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25812;

architecture SYN_ARCHBEH of nd2_25812 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25811 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25811;

architecture SYN_ARCHBEH of nd2_25811 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25810 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25810;

architecture SYN_ARCHBEH of nd2_25810 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25809 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25809;

architecture SYN_ARCHBEH of nd2_25809 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25808 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25808;

architecture SYN_ARCHBEH of nd2_25808 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25807 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25807;

architecture SYN_ARCHBEH of nd2_25807 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25806 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25806;

architecture SYN_ARCHBEH of nd2_25806 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25805 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25805;

architecture SYN_ARCHBEH of nd2_25805 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25804 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25804;

architecture SYN_ARCHBEH of nd2_25804 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25803 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25803;

architecture SYN_ARCHBEH of nd2_25803 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25802 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25802;

architecture SYN_ARCHBEH of nd2_25802 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25801 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25801;

architecture SYN_ARCHBEH of nd2_25801 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25800 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25800;

architecture SYN_ARCHBEH of nd2_25800 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25799 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25799;

architecture SYN_ARCHBEH of nd2_25799 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25798 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25798;

architecture SYN_ARCHBEH of nd2_25798 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25797 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25797;

architecture SYN_ARCHBEH of nd2_25797 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25796 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25796;

architecture SYN_ARCHBEH of nd2_25796 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25795 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25795;

architecture SYN_ARCHBEH of nd2_25795 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25794 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25794;

architecture SYN_ARCHBEH of nd2_25794 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25793 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25793;

architecture SYN_ARCHBEH of nd2_25793 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25792 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25792;

architecture SYN_ARCHBEH of nd2_25792 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25791 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25791;

architecture SYN_ARCHBEH of nd2_25791 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25790 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25790;

architecture SYN_ARCHBEH of nd2_25790 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25789 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25789;

architecture SYN_ARCHBEH of nd2_25789 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25788 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25788;

architecture SYN_ARCHBEH of nd2_25788 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25787 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25787;

architecture SYN_ARCHBEH of nd2_25787 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25786 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25786;

architecture SYN_ARCHBEH of nd2_25786 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25785 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25785;

architecture SYN_ARCHBEH of nd2_25785 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25784 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25784;

architecture SYN_ARCHBEH of nd2_25784 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25783 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25783;

architecture SYN_ARCHBEH of nd2_25783 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25782 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25782;

architecture SYN_ARCHBEH of nd2_25782 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25781 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25781;

architecture SYN_ARCHBEH of nd2_25781 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25780 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25780;

architecture SYN_ARCHBEH of nd2_25780 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25779 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25779;

architecture SYN_ARCHBEH of nd2_25779 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25778 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25778;

architecture SYN_ARCHBEH of nd2_25778 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25777 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25777;

architecture SYN_ARCHBEH of nd2_25777 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25776 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25776;

architecture SYN_ARCHBEH of nd2_25776 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25775 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25775;

architecture SYN_ARCHBEH of nd2_25775 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25774 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25774;

architecture SYN_ARCHBEH of nd2_25774 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25773 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25773;

architecture SYN_ARCHBEH of nd2_25773 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25772 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25772;

architecture SYN_ARCHBEH of nd2_25772 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25771 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25771;

architecture SYN_ARCHBEH of nd2_25771 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25770 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25770;

architecture SYN_ARCHBEH of nd2_25770 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25769 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25769;

architecture SYN_ARCHBEH of nd2_25769 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25768 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25768;

architecture SYN_ARCHBEH of nd2_25768 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25767 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25767;

architecture SYN_ARCHBEH of nd2_25767 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25766 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25766;

architecture SYN_ARCHBEH of nd2_25766 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25765 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25765;

architecture SYN_ARCHBEH of nd2_25765 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25764 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25764;

architecture SYN_ARCHBEH of nd2_25764 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25763 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25763;

architecture SYN_ARCHBEH of nd2_25763 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25762 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25762;

architecture SYN_ARCHBEH of nd2_25762 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25761 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25761;

architecture SYN_ARCHBEH of nd2_25761 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25760 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25760;

architecture SYN_ARCHBEH of nd2_25760 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25759 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25759;

architecture SYN_ARCHBEH of nd2_25759 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25758 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25758;

architecture SYN_ARCHBEH of nd2_25758 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25757 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25757;

architecture SYN_ARCHBEH of nd2_25757 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25756 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25756;

architecture SYN_ARCHBEH of nd2_25756 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25755 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25755;

architecture SYN_ARCHBEH of nd2_25755 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25754 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25754;

architecture SYN_ARCHBEH of nd2_25754 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25753 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25753;

architecture SYN_ARCHBEH of nd2_25753 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25752 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25752;

architecture SYN_ARCHBEH of nd2_25752 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25751 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25751;

architecture SYN_ARCHBEH of nd2_25751 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25750 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25750;

architecture SYN_ARCHBEH of nd2_25750 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25749 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25749;

architecture SYN_ARCHBEH of nd2_25749 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25748 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25748;

architecture SYN_ARCHBEH of nd2_25748 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25747 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25747;

architecture SYN_ARCHBEH of nd2_25747 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25746 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25746;

architecture SYN_ARCHBEH of nd2_25746 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25745 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25745;

architecture SYN_ARCHBEH of nd2_25745 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25744 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25744;

architecture SYN_ARCHBEH of nd2_25744 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25743 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25743;

architecture SYN_ARCHBEH of nd2_25743 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25742 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25742;

architecture SYN_ARCHBEH of nd2_25742 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25741 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25741;

architecture SYN_ARCHBEH of nd2_25741 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25740 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25740;

architecture SYN_ARCHBEH of nd2_25740 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25739 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25739;

architecture SYN_ARCHBEH of nd2_25739 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25738 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25738;

architecture SYN_ARCHBEH of nd2_25738 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25737 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25737;

architecture SYN_ARCHBEH of nd2_25737 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25736 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25736;

architecture SYN_ARCHBEH of nd2_25736 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25735 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25735;

architecture SYN_ARCHBEH of nd2_25735 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25734 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25734;

architecture SYN_ARCHBEH of nd2_25734 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25733 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25733;

architecture SYN_ARCHBEH of nd2_25733 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25732 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25732;

architecture SYN_ARCHBEH of nd2_25732 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25731 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25731;

architecture SYN_ARCHBEH of nd2_25731 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25730 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25730;

architecture SYN_ARCHBEH of nd2_25730 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25729 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25729;

architecture SYN_ARCHBEH of nd2_25729 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25728 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25728;

architecture SYN_ARCHBEH of nd2_25728 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25727 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25727;

architecture SYN_ARCHBEH of nd2_25727 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25726 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25726;

architecture SYN_ARCHBEH of nd2_25726 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25725 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25725;

architecture SYN_ARCHBEH of nd2_25725 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25724 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25724;

architecture SYN_ARCHBEH of nd2_25724 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25723 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25723;

architecture SYN_ARCHBEH of nd2_25723 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25722 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25722;

architecture SYN_ARCHBEH of nd2_25722 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25721 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25721;

architecture SYN_ARCHBEH of nd2_25721 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25720 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25720;

architecture SYN_ARCHBEH of nd2_25720 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25719 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25719;

architecture SYN_ARCHBEH of nd2_25719 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25718 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25718;

architecture SYN_ARCHBEH of nd2_25718 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25717 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25717;

architecture SYN_ARCHBEH of nd2_25717 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25716 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25716;

architecture SYN_ARCHBEH of nd2_25716 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25715 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25715;

architecture SYN_ARCHBEH of nd2_25715 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25714 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25714;

architecture SYN_ARCHBEH of nd2_25714 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25713 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25713;

architecture SYN_ARCHBEH of nd2_25713 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25712 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25712;

architecture SYN_ARCHBEH of nd2_25712 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25711 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25711;

architecture SYN_ARCHBEH of nd2_25711 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25710 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25710;

architecture SYN_ARCHBEH of nd2_25710 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25709 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25709;

architecture SYN_ARCHBEH of nd2_25709 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25708 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25708;

architecture SYN_ARCHBEH of nd2_25708 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25707 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25707;

architecture SYN_ARCHBEH of nd2_25707 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25706 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25706;

architecture SYN_ARCHBEH of nd2_25706 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25705 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25705;

architecture SYN_ARCHBEH of nd2_25705 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25704 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25704;

architecture SYN_ARCHBEH of nd2_25704 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25703 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25703;

architecture SYN_ARCHBEH of nd2_25703 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25702 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25702;

architecture SYN_ARCHBEH of nd2_25702 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25701 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25701;

architecture SYN_ARCHBEH of nd2_25701 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25700 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25700;

architecture SYN_ARCHBEH of nd2_25700 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25699 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25699;

architecture SYN_ARCHBEH of nd2_25699 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25698 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25698;

architecture SYN_ARCHBEH of nd2_25698 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25697 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25697;

architecture SYN_ARCHBEH of nd2_25697 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25696 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25696;

architecture SYN_ARCHBEH of nd2_25696 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25695 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25695;

architecture SYN_ARCHBEH of nd2_25695 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25694 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25694;

architecture SYN_ARCHBEH of nd2_25694 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25693 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25693;

architecture SYN_ARCHBEH of nd2_25693 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25692 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25692;

architecture SYN_ARCHBEH of nd2_25692 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25691 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25691;

architecture SYN_ARCHBEH of nd2_25691 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25690 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25690;

architecture SYN_ARCHBEH of nd2_25690 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25689 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25689;

architecture SYN_ARCHBEH of nd2_25689 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25688 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25688;

architecture SYN_ARCHBEH of nd2_25688 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25687 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25687;

architecture SYN_ARCHBEH of nd2_25687 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25686 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25686;

architecture SYN_ARCHBEH of nd2_25686 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25685 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25685;

architecture SYN_ARCHBEH of nd2_25685 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25684 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25684;

architecture SYN_ARCHBEH of nd2_25684 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25683 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25683;

architecture SYN_ARCHBEH of nd2_25683 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25682 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25682;

architecture SYN_ARCHBEH of nd2_25682 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25681 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25681;

architecture SYN_ARCHBEH of nd2_25681 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25680 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25680;

architecture SYN_ARCHBEH of nd2_25680 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25679 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25679;

architecture SYN_ARCHBEH of nd2_25679 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25678 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25678;

architecture SYN_ARCHBEH of nd2_25678 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25677 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25677;

architecture SYN_ARCHBEH of nd2_25677 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25676 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25676;

architecture SYN_ARCHBEH of nd2_25676 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25675 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25675;

architecture SYN_ARCHBEH of nd2_25675 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25674 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25674;

architecture SYN_ARCHBEH of nd2_25674 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25673 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25673;

architecture SYN_ARCHBEH of nd2_25673 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25672 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25672;

architecture SYN_ARCHBEH of nd2_25672 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25671 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25671;

architecture SYN_ARCHBEH of nd2_25671 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25670 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25670;

architecture SYN_ARCHBEH of nd2_25670 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25669 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25669;

architecture SYN_ARCHBEH of nd2_25669 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25668 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25668;

architecture SYN_ARCHBEH of nd2_25668 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25667 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25667;

architecture SYN_ARCHBEH of nd2_25667 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25666 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25666;

architecture SYN_ARCHBEH of nd2_25666 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25665 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25665;

architecture SYN_ARCHBEH of nd2_25665 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25664 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25664;

architecture SYN_ARCHBEH of nd2_25664 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25663 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25663;

architecture SYN_ARCHBEH of nd2_25663 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25662 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25662;

architecture SYN_ARCHBEH of nd2_25662 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25661 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25661;

architecture SYN_ARCHBEH of nd2_25661 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25660 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25660;

architecture SYN_ARCHBEH of nd2_25660 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25659 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25659;

architecture SYN_ARCHBEH of nd2_25659 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25658 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25658;

architecture SYN_ARCHBEH of nd2_25658 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25657 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25657;

architecture SYN_ARCHBEH of nd2_25657 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25656 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25656;

architecture SYN_ARCHBEH of nd2_25656 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25655 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25655;

architecture SYN_ARCHBEH of nd2_25655 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25654 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25654;

architecture SYN_ARCHBEH of nd2_25654 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25653 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25653;

architecture SYN_ARCHBEH of nd2_25653 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25652 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25652;

architecture SYN_ARCHBEH of nd2_25652 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25651 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25651;

architecture SYN_ARCHBEH of nd2_25651 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25650 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25650;

architecture SYN_ARCHBEH of nd2_25650 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25649 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25649;

architecture SYN_ARCHBEH of nd2_25649 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25648 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25648;

architecture SYN_ARCHBEH of nd2_25648 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25647 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25647;

architecture SYN_ARCHBEH of nd2_25647 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25646 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25646;

architecture SYN_ARCHBEH of nd2_25646 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25645 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25645;

architecture SYN_ARCHBEH of nd2_25645 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25644 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25644;

architecture SYN_ARCHBEH of nd2_25644 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25643 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25643;

architecture SYN_ARCHBEH of nd2_25643 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25642 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25642;

architecture SYN_ARCHBEH of nd2_25642 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25641 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25641;

architecture SYN_ARCHBEH of nd2_25641 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25640 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25640;

architecture SYN_ARCHBEH of nd2_25640 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25639 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25639;

architecture SYN_ARCHBEH of nd2_25639 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25638 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25638;

architecture SYN_ARCHBEH of nd2_25638 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25637 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25637;

architecture SYN_ARCHBEH of nd2_25637 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25636 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25636;

architecture SYN_ARCHBEH of nd2_25636 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25635 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25635;

architecture SYN_ARCHBEH of nd2_25635 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25634 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25634;

architecture SYN_ARCHBEH of nd2_25634 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25633 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25633;

architecture SYN_ARCHBEH of nd2_25633 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25632 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25632;

architecture SYN_ARCHBEH of nd2_25632 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25631 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25631;

architecture SYN_ARCHBEH of nd2_25631 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25630 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25630;

architecture SYN_ARCHBEH of nd2_25630 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25629 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25629;

architecture SYN_ARCHBEH of nd2_25629 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25628 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25628;

architecture SYN_ARCHBEH of nd2_25628 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25627 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25627;

architecture SYN_ARCHBEH of nd2_25627 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25626 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25626;

architecture SYN_ARCHBEH of nd2_25626 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25625 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25625;

architecture SYN_ARCHBEH of nd2_25625 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25624 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25624;

architecture SYN_ARCHBEH of nd2_25624 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25623 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25623;

architecture SYN_ARCHBEH of nd2_25623 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25622 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25622;

architecture SYN_ARCHBEH of nd2_25622 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25621 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25621;

architecture SYN_ARCHBEH of nd2_25621 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25620 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25620;

architecture SYN_ARCHBEH of nd2_25620 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25619 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25619;

architecture SYN_ARCHBEH of nd2_25619 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25618 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25618;

architecture SYN_ARCHBEH of nd2_25618 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25617 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25617;

architecture SYN_ARCHBEH of nd2_25617 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25616 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25616;

architecture SYN_ARCHBEH of nd2_25616 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25615 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25615;

architecture SYN_ARCHBEH of nd2_25615 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25614 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25614;

architecture SYN_ARCHBEH of nd2_25614 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25613 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25613;

architecture SYN_ARCHBEH of nd2_25613 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25612 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25612;

architecture SYN_ARCHBEH of nd2_25612 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25611 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25611;

architecture SYN_ARCHBEH of nd2_25611 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25610 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25610;

architecture SYN_ARCHBEH of nd2_25610 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25609 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25609;

architecture SYN_ARCHBEH of nd2_25609 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25608 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25608;

architecture SYN_ARCHBEH of nd2_25608 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25607 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25607;

architecture SYN_ARCHBEH of nd2_25607 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25606 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25606;

architecture SYN_ARCHBEH of nd2_25606 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25605 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25605;

architecture SYN_ARCHBEH of nd2_25605 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25604 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25604;

architecture SYN_ARCHBEH of nd2_25604 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25603 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25603;

architecture SYN_ARCHBEH of nd2_25603 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25602 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25602;

architecture SYN_ARCHBEH of nd2_25602 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25601 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25601;

architecture SYN_ARCHBEH of nd2_25601 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25600 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25600;

architecture SYN_ARCHBEH of nd2_25600 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25599 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25599;

architecture SYN_ARCHBEH of nd2_25599 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25598 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25598;

architecture SYN_ARCHBEH of nd2_25598 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25597 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25597;

architecture SYN_ARCHBEH of nd2_25597 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25596 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25596;

architecture SYN_ARCHBEH of nd2_25596 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25595 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25595;

architecture SYN_ARCHBEH of nd2_25595 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25594 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25594;

architecture SYN_ARCHBEH of nd2_25594 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25593 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25593;

architecture SYN_ARCHBEH of nd2_25593 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25592 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25592;

architecture SYN_ARCHBEH of nd2_25592 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25591 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25591;

architecture SYN_ARCHBEH of nd2_25591 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25590 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25590;

architecture SYN_ARCHBEH of nd2_25590 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25589 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25589;

architecture SYN_ARCHBEH of nd2_25589 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25588 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25588;

architecture SYN_ARCHBEH of nd2_25588 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25587 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25587;

architecture SYN_ARCHBEH of nd2_25587 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25586 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25586;

architecture SYN_ARCHBEH of nd2_25586 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25585 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25585;

architecture SYN_ARCHBEH of nd2_25585 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25584 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25584;

architecture SYN_ARCHBEH of nd2_25584 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25583 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25583;

architecture SYN_ARCHBEH of nd2_25583 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25582 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25582;

architecture SYN_ARCHBEH of nd2_25582 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25581 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25581;

architecture SYN_ARCHBEH of nd2_25581 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25580 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25580;

architecture SYN_ARCHBEH of nd2_25580 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25579 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25579;

architecture SYN_ARCHBEH of nd2_25579 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25578 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25578;

architecture SYN_ARCHBEH of nd2_25578 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25577 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25577;

architecture SYN_ARCHBEH of nd2_25577 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25576 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25576;

architecture SYN_ARCHBEH of nd2_25576 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25575 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25575;

architecture SYN_ARCHBEH of nd2_25575 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25574 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25574;

architecture SYN_ARCHBEH of nd2_25574 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25573 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25573;

architecture SYN_ARCHBEH of nd2_25573 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25572 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25572;

architecture SYN_ARCHBEH of nd2_25572 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25571 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25571;

architecture SYN_ARCHBEH of nd2_25571 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25570 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25570;

architecture SYN_ARCHBEH of nd2_25570 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25569 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25569;

architecture SYN_ARCHBEH of nd2_25569 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25568 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25568;

architecture SYN_ARCHBEH of nd2_25568 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25567 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25567;

architecture SYN_ARCHBEH of nd2_25567 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25566 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25566;

architecture SYN_ARCHBEH of nd2_25566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25565 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25565;

architecture SYN_ARCHBEH of nd2_25565 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25564 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25564;

architecture SYN_ARCHBEH of nd2_25564 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25563 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25563;

architecture SYN_ARCHBEH of nd2_25563 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25562 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25562;

architecture SYN_ARCHBEH of nd2_25562 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25561 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25561;

architecture SYN_ARCHBEH of nd2_25561 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25560 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25560;

architecture SYN_ARCHBEH of nd2_25560 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25559 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25559;

architecture SYN_ARCHBEH of nd2_25559 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25558 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25558;

architecture SYN_ARCHBEH of nd2_25558 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25557 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25557;

architecture SYN_ARCHBEH of nd2_25557 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25556 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25556;

architecture SYN_ARCHBEH of nd2_25556 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25555 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25555;

architecture SYN_ARCHBEH of nd2_25555 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25554 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25554;

architecture SYN_ARCHBEH of nd2_25554 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25553 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25553;

architecture SYN_ARCHBEH of nd2_25553 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25552 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25552;

architecture SYN_ARCHBEH of nd2_25552 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25551 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25551;

architecture SYN_ARCHBEH of nd2_25551 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25550 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25550;

architecture SYN_ARCHBEH of nd2_25550 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25549 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25549;

architecture SYN_ARCHBEH of nd2_25549 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25548 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25548;

architecture SYN_ARCHBEH of nd2_25548 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25547 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25547;

architecture SYN_ARCHBEH of nd2_25547 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25546 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25546;

architecture SYN_ARCHBEH of nd2_25546 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25545 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25545;

architecture SYN_ARCHBEH of nd2_25545 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25544 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25544;

architecture SYN_ARCHBEH of nd2_25544 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25543 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25543;

architecture SYN_ARCHBEH of nd2_25543 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25542 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25542;

architecture SYN_ARCHBEH of nd2_25542 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25541 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25541;

architecture SYN_ARCHBEH of nd2_25541 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25540 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25540;

architecture SYN_ARCHBEH of nd2_25540 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25539 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25539;

architecture SYN_ARCHBEH of nd2_25539 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25538 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25538;

architecture SYN_ARCHBEH of nd2_25538 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25537 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25537;

architecture SYN_ARCHBEH of nd2_25537 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25536 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25536;

architecture SYN_ARCHBEH of nd2_25536 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25535 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25535;

architecture SYN_ARCHBEH of nd2_25535 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25534 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25534;

architecture SYN_ARCHBEH of nd2_25534 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25533 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25533;

architecture SYN_ARCHBEH of nd2_25533 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25532 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25532;

architecture SYN_ARCHBEH of nd2_25532 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25531 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25531;

architecture SYN_ARCHBEH of nd2_25531 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25530 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25530;

architecture SYN_ARCHBEH of nd2_25530 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25529 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25529;

architecture SYN_ARCHBEH of nd2_25529 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25528 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25528;

architecture SYN_ARCHBEH of nd2_25528 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25527 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25527;

architecture SYN_ARCHBEH of nd2_25527 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25526 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25526;

architecture SYN_ARCHBEH of nd2_25526 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25525 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25525;

architecture SYN_ARCHBEH of nd2_25525 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25524 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25524;

architecture SYN_ARCHBEH of nd2_25524 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25523 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25523;

architecture SYN_ARCHBEH of nd2_25523 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25522 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25522;

architecture SYN_ARCHBEH of nd2_25522 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25521 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25521;

architecture SYN_ARCHBEH of nd2_25521 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25520 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25520;

architecture SYN_ARCHBEH of nd2_25520 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25519 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25519;

architecture SYN_ARCHBEH of nd2_25519 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25518 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25518;

architecture SYN_ARCHBEH of nd2_25518 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25517 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25517;

architecture SYN_ARCHBEH of nd2_25517 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25516 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25516;

architecture SYN_ARCHBEH of nd2_25516 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25515 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25515;

architecture SYN_ARCHBEH of nd2_25515 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25514 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25514;

architecture SYN_ARCHBEH of nd2_25514 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25513 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25513;

architecture SYN_ARCHBEH of nd2_25513 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25512 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25512;

architecture SYN_ARCHBEH of nd2_25512 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25511 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25511;

architecture SYN_ARCHBEH of nd2_25511 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25510 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25510;

architecture SYN_ARCHBEH of nd2_25510 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25509 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25509;

architecture SYN_ARCHBEH of nd2_25509 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25508 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25508;

architecture SYN_ARCHBEH of nd2_25508 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25507 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25507;

architecture SYN_ARCHBEH of nd2_25507 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25506 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25506;

architecture SYN_ARCHBEH of nd2_25506 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25505 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25505;

architecture SYN_ARCHBEH of nd2_25505 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25504 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25504;

architecture SYN_ARCHBEH of nd2_25504 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25503 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25503;

architecture SYN_ARCHBEH of nd2_25503 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25502 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25502;

architecture SYN_ARCHBEH of nd2_25502 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25501 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25501;

architecture SYN_ARCHBEH of nd2_25501 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25500 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25500;

architecture SYN_ARCHBEH of nd2_25500 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25499 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25499;

architecture SYN_ARCHBEH of nd2_25499 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25498 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25498;

architecture SYN_ARCHBEH of nd2_25498 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25497 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25497;

architecture SYN_ARCHBEH of nd2_25497 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25496 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25496;

architecture SYN_ARCHBEH of nd2_25496 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25495 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25495;

architecture SYN_ARCHBEH of nd2_25495 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25494 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25494;

architecture SYN_ARCHBEH of nd2_25494 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25493 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25493;

architecture SYN_ARCHBEH of nd2_25493 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25492 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25492;

architecture SYN_ARCHBEH of nd2_25492 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25491 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25491;

architecture SYN_ARCHBEH of nd2_25491 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25490 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25490;

architecture SYN_ARCHBEH of nd2_25490 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25489 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25489;

architecture SYN_ARCHBEH of nd2_25489 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25488 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25488;

architecture SYN_ARCHBEH of nd2_25488 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25487 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25487;

architecture SYN_ARCHBEH of nd2_25487 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25486 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25486;

architecture SYN_ARCHBEH of nd2_25486 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25485 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25485;

architecture SYN_ARCHBEH of nd2_25485 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25484 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25484;

architecture SYN_ARCHBEH of nd2_25484 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25483 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25483;

architecture SYN_ARCHBEH of nd2_25483 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25482 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25482;

architecture SYN_ARCHBEH of nd2_25482 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25481 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25481;

architecture SYN_ARCHBEH of nd2_25481 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25480 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25480;

architecture SYN_ARCHBEH of nd2_25480 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25479 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25479;

architecture SYN_ARCHBEH of nd2_25479 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25478 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25478;

architecture SYN_ARCHBEH of nd2_25478 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25477 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25477;

architecture SYN_ARCHBEH of nd2_25477 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25476 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25476;

architecture SYN_ARCHBEH of nd2_25476 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25475 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25475;

architecture SYN_ARCHBEH of nd2_25475 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25474 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25474;

architecture SYN_ARCHBEH of nd2_25474 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25473 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25473;

architecture SYN_ARCHBEH of nd2_25473 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25472 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25472;

architecture SYN_ARCHBEH of nd2_25472 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25471 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25471;

architecture SYN_ARCHBEH of nd2_25471 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25470 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25470;

architecture SYN_ARCHBEH of nd2_25470 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25469 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25469;

architecture SYN_ARCHBEH of nd2_25469 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25468 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25468;

architecture SYN_ARCHBEH of nd2_25468 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25467 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25467;

architecture SYN_ARCHBEH of nd2_25467 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25466 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25466;

architecture SYN_ARCHBEH of nd2_25466 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25465 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25465;

architecture SYN_ARCHBEH of nd2_25465 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25464 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25464;

architecture SYN_ARCHBEH of nd2_25464 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25463 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25463;

architecture SYN_ARCHBEH of nd2_25463 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25462 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25462;

architecture SYN_ARCHBEH of nd2_25462 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25461 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25461;

architecture SYN_ARCHBEH of nd2_25461 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25460 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25460;

architecture SYN_ARCHBEH of nd2_25460 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25459 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25459;

architecture SYN_ARCHBEH of nd2_25459 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25458 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25458;

architecture SYN_ARCHBEH of nd2_25458 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25457 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25457;

architecture SYN_ARCHBEH of nd2_25457 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25456 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25456;

architecture SYN_ARCHBEH of nd2_25456 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25455 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25455;

architecture SYN_ARCHBEH of nd2_25455 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25454 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25454;

architecture SYN_ARCHBEH of nd2_25454 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25453 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25453;

architecture SYN_ARCHBEH of nd2_25453 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25452 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25452;

architecture SYN_ARCHBEH of nd2_25452 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25451 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25451;

architecture SYN_ARCHBEH of nd2_25451 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25450 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25450;

architecture SYN_ARCHBEH of nd2_25450 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25449 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25449;

architecture SYN_ARCHBEH of nd2_25449 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25448 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25448;

architecture SYN_ARCHBEH of nd2_25448 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25447 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25447;

architecture SYN_ARCHBEH of nd2_25447 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25446 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25446;

architecture SYN_ARCHBEH of nd2_25446 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25445 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25445;

architecture SYN_ARCHBEH of nd2_25445 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25444 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25444;

architecture SYN_ARCHBEH of nd2_25444 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25443 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25443;

architecture SYN_ARCHBEH of nd2_25443 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25442 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25442;

architecture SYN_ARCHBEH of nd2_25442 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25441 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25441;

architecture SYN_ARCHBEH of nd2_25441 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25440 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25440;

architecture SYN_ARCHBEH of nd2_25440 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25439 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25439;

architecture SYN_ARCHBEH of nd2_25439 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25438 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25438;

architecture SYN_ARCHBEH of nd2_25438 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25437 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25437;

architecture SYN_ARCHBEH of nd2_25437 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25436 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25436;

architecture SYN_ARCHBEH of nd2_25436 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25435 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25435;

architecture SYN_ARCHBEH of nd2_25435 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25434 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25434;

architecture SYN_ARCHBEH of nd2_25434 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25433 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25433;

architecture SYN_ARCHBEH of nd2_25433 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25432 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25432;

architecture SYN_ARCHBEH of nd2_25432 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25431 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25431;

architecture SYN_ARCHBEH of nd2_25431 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25430 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25430;

architecture SYN_ARCHBEH of nd2_25430 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25429 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25429;

architecture SYN_ARCHBEH of nd2_25429 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25428 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25428;

architecture SYN_ARCHBEH of nd2_25428 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25427 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25427;

architecture SYN_ARCHBEH of nd2_25427 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25426 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25426;

architecture SYN_ARCHBEH of nd2_25426 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25425 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25425;

architecture SYN_ARCHBEH of nd2_25425 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25424 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25424;

architecture SYN_ARCHBEH of nd2_25424 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25423 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25423;

architecture SYN_ARCHBEH of nd2_25423 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25422 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25422;

architecture SYN_ARCHBEH of nd2_25422 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25421 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25421;

architecture SYN_ARCHBEH of nd2_25421 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25420 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25420;

architecture SYN_ARCHBEH of nd2_25420 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25419 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25419;

architecture SYN_ARCHBEH of nd2_25419 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25418 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25418;

architecture SYN_ARCHBEH of nd2_25418 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25417 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25417;

architecture SYN_ARCHBEH of nd2_25417 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25416 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25416;

architecture SYN_ARCHBEH of nd2_25416 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25415 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25415;

architecture SYN_ARCHBEH of nd2_25415 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25414 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25414;

architecture SYN_ARCHBEH of nd2_25414 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25413 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25413;

architecture SYN_ARCHBEH of nd2_25413 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25412 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25412;

architecture SYN_ARCHBEH of nd2_25412 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25411 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25411;

architecture SYN_ARCHBEH of nd2_25411 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25410 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25410;

architecture SYN_ARCHBEH of nd2_25410 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25409 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25409;

architecture SYN_ARCHBEH of nd2_25409 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25408 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25408;

architecture SYN_ARCHBEH of nd2_25408 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25407 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25407;

architecture SYN_ARCHBEH of nd2_25407 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25406 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25406;

architecture SYN_ARCHBEH of nd2_25406 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25405 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25405;

architecture SYN_ARCHBEH of nd2_25405 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25404 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25404;

architecture SYN_ARCHBEH of nd2_25404 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25403 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25403;

architecture SYN_ARCHBEH of nd2_25403 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25402 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25402;

architecture SYN_ARCHBEH of nd2_25402 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25401 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25401;

architecture SYN_ARCHBEH of nd2_25401 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25400 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25400;

architecture SYN_ARCHBEH of nd2_25400 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25399 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25399;

architecture SYN_ARCHBEH of nd2_25399 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25398 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25398;

architecture SYN_ARCHBEH of nd2_25398 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25397 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25397;

architecture SYN_ARCHBEH of nd2_25397 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25396 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25396;

architecture SYN_ARCHBEH of nd2_25396 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25395 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25395;

architecture SYN_ARCHBEH of nd2_25395 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25394 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25394;

architecture SYN_ARCHBEH of nd2_25394 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25393 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25393;

architecture SYN_ARCHBEH of nd2_25393 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25392 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25392;

architecture SYN_ARCHBEH of nd2_25392 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25391 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25391;

architecture SYN_ARCHBEH of nd2_25391 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25390 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25390;

architecture SYN_ARCHBEH of nd2_25390 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25389 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25389;

architecture SYN_ARCHBEH of nd2_25389 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25388 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25388;

architecture SYN_ARCHBEH of nd2_25388 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25387 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25387;

architecture SYN_ARCHBEH of nd2_25387 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25386 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25386;

architecture SYN_ARCHBEH of nd2_25386 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25385 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25385;

architecture SYN_ARCHBEH of nd2_25385 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25384 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25384;

architecture SYN_ARCHBEH of nd2_25384 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25383 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25383;

architecture SYN_ARCHBEH of nd2_25383 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25382 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25382;

architecture SYN_ARCHBEH of nd2_25382 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25381 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25381;

architecture SYN_ARCHBEH of nd2_25381 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25380 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25380;

architecture SYN_ARCHBEH of nd2_25380 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25379 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25379;

architecture SYN_ARCHBEH of nd2_25379 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25378 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25378;

architecture SYN_ARCHBEH of nd2_25378 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25377 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25377;

architecture SYN_ARCHBEH of nd2_25377 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25376 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25376;

architecture SYN_ARCHBEH of nd2_25376 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25375 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25375;

architecture SYN_ARCHBEH of nd2_25375 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25374 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25374;

architecture SYN_ARCHBEH of nd2_25374 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25373 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25373;

architecture SYN_ARCHBEH of nd2_25373 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25372 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25372;

architecture SYN_ARCHBEH of nd2_25372 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25371 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25371;

architecture SYN_ARCHBEH of nd2_25371 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25370 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25370;

architecture SYN_ARCHBEH of nd2_25370 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25369 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25369;

architecture SYN_ARCHBEH of nd2_25369 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25368 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25368;

architecture SYN_ARCHBEH of nd2_25368 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25367 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25367;

architecture SYN_ARCHBEH of nd2_25367 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25366 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25366;

architecture SYN_ARCHBEH of nd2_25366 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25365 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25365;

architecture SYN_ARCHBEH of nd2_25365 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25364 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25364;

architecture SYN_ARCHBEH of nd2_25364 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25363 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25363;

architecture SYN_ARCHBEH of nd2_25363 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25362 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25362;

architecture SYN_ARCHBEH of nd2_25362 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25361 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25361;

architecture SYN_ARCHBEH of nd2_25361 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25360 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25360;

architecture SYN_ARCHBEH of nd2_25360 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25359 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25359;

architecture SYN_ARCHBEH of nd2_25359 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25358 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25358;

architecture SYN_ARCHBEH of nd2_25358 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25357 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25357;

architecture SYN_ARCHBEH of nd2_25357 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25356 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25356;

architecture SYN_ARCHBEH of nd2_25356 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25355 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25355;

architecture SYN_ARCHBEH of nd2_25355 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25354 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25354;

architecture SYN_ARCHBEH of nd2_25354 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25353 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25353;

architecture SYN_ARCHBEH of nd2_25353 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25352 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25352;

architecture SYN_ARCHBEH of nd2_25352 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25351 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25351;

architecture SYN_ARCHBEH of nd2_25351 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25350 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25350;

architecture SYN_ARCHBEH of nd2_25350 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25349 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25349;

architecture SYN_ARCHBEH of nd2_25349 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25348 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25348;

architecture SYN_ARCHBEH of nd2_25348 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25347 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25347;

architecture SYN_ARCHBEH of nd2_25347 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25346 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25346;

architecture SYN_ARCHBEH of nd2_25346 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25345 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25345;

architecture SYN_ARCHBEH of nd2_25345 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25344 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25344;

architecture SYN_ARCHBEH of nd2_25344 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25343 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25343;

architecture SYN_ARCHBEH of nd2_25343 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25342 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25342;

architecture SYN_ARCHBEH of nd2_25342 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25341 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25341;

architecture SYN_ARCHBEH of nd2_25341 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25340 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25340;

architecture SYN_ARCHBEH of nd2_25340 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25339 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25339;

architecture SYN_ARCHBEH of nd2_25339 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25338 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25338;

architecture SYN_ARCHBEH of nd2_25338 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25337 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25337;

architecture SYN_ARCHBEH of nd2_25337 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25336 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25336;

architecture SYN_ARCHBEH of nd2_25336 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25335 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25335;

architecture SYN_ARCHBEH of nd2_25335 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25334 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25334;

architecture SYN_ARCHBEH of nd2_25334 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25333 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25333;

architecture SYN_ARCHBEH of nd2_25333 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25332 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25332;

architecture SYN_ARCHBEH of nd2_25332 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25331 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25331;

architecture SYN_ARCHBEH of nd2_25331 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25330 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25330;

architecture SYN_ARCHBEH of nd2_25330 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25329 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25329;

architecture SYN_ARCHBEH of nd2_25329 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25328 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25328;

architecture SYN_ARCHBEH of nd2_25328 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25327 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25327;

architecture SYN_ARCHBEH of nd2_25327 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25326 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25326;

architecture SYN_ARCHBEH of nd2_25326 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25325 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25325;

architecture SYN_ARCHBEH of nd2_25325 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25324 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25324;

architecture SYN_ARCHBEH of nd2_25324 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25323 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25323;

architecture SYN_ARCHBEH of nd2_25323 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25322 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25322;

architecture SYN_ARCHBEH of nd2_25322 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25321 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25321;

architecture SYN_ARCHBEH of nd2_25321 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25320 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25320;

architecture SYN_ARCHBEH of nd2_25320 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25319 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25319;

architecture SYN_ARCHBEH of nd2_25319 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25318 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25318;

architecture SYN_ARCHBEH of nd2_25318 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25317 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25317;

architecture SYN_ARCHBEH of nd2_25317 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25316 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25316;

architecture SYN_ARCHBEH of nd2_25316 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25315 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25315;

architecture SYN_ARCHBEH of nd2_25315 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25314 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25314;

architecture SYN_ARCHBEH of nd2_25314 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25313 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25313;

architecture SYN_ARCHBEH of nd2_25313 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25312 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25312;

architecture SYN_ARCHBEH of nd2_25312 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25311 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25311;

architecture SYN_ARCHBEH of nd2_25311 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25310 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25310;

architecture SYN_ARCHBEH of nd2_25310 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25309 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25309;

architecture SYN_ARCHBEH of nd2_25309 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25308 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25308;

architecture SYN_ARCHBEH of nd2_25308 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25307 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25307;

architecture SYN_ARCHBEH of nd2_25307 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25306 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25306;

architecture SYN_ARCHBEH of nd2_25306 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25305 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25305;

architecture SYN_ARCHBEH of nd2_25305 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25304 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25304;

architecture SYN_ARCHBEH of nd2_25304 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25303 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25303;

architecture SYN_ARCHBEH of nd2_25303 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25302 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25302;

architecture SYN_ARCHBEH of nd2_25302 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25301 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25301;

architecture SYN_ARCHBEH of nd2_25301 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25300 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25300;

architecture SYN_ARCHBEH of nd2_25300 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25299 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25299;

architecture SYN_ARCHBEH of nd2_25299 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25298 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25298;

architecture SYN_ARCHBEH of nd2_25298 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25297 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25297;

architecture SYN_ARCHBEH of nd2_25297 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25296 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25296;

architecture SYN_ARCHBEH of nd2_25296 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25295 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25295;

architecture SYN_ARCHBEH of nd2_25295 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25294 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25294;

architecture SYN_ARCHBEH of nd2_25294 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25293 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25293;

architecture SYN_ARCHBEH of nd2_25293 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25292 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25292;

architecture SYN_ARCHBEH of nd2_25292 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25291 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25291;

architecture SYN_ARCHBEH of nd2_25291 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25290 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25290;

architecture SYN_ARCHBEH of nd2_25290 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25289 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25289;

architecture SYN_ARCHBEH of nd2_25289 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25288 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25288;

architecture SYN_ARCHBEH of nd2_25288 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25287 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25287;

architecture SYN_ARCHBEH of nd2_25287 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25286 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25286;

architecture SYN_ARCHBEH of nd2_25286 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25285 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25285;

architecture SYN_ARCHBEH of nd2_25285 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25284 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25284;

architecture SYN_ARCHBEH of nd2_25284 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25283 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25283;

architecture SYN_ARCHBEH of nd2_25283 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25282 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25282;

architecture SYN_ARCHBEH of nd2_25282 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25281 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25281;

architecture SYN_ARCHBEH of nd2_25281 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25280 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25280;

architecture SYN_ARCHBEH of nd2_25280 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25279 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25279;

architecture SYN_ARCHBEH of nd2_25279 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25278 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25278;

architecture SYN_ARCHBEH of nd2_25278 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25277 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25277;

architecture SYN_ARCHBEH of nd2_25277 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25276 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25276;

architecture SYN_ARCHBEH of nd2_25276 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25275 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25275;

architecture SYN_ARCHBEH of nd2_25275 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25274 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25274;

architecture SYN_ARCHBEH of nd2_25274 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25273 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25273;

architecture SYN_ARCHBEH of nd2_25273 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25272 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25272;

architecture SYN_ARCHBEH of nd2_25272 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25271 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25271;

architecture SYN_ARCHBEH of nd2_25271 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25270 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25270;

architecture SYN_ARCHBEH of nd2_25270 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25269 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25269;

architecture SYN_ARCHBEH of nd2_25269 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25268 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25268;

architecture SYN_ARCHBEH of nd2_25268 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25267 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25267;

architecture SYN_ARCHBEH of nd2_25267 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25266 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25266;

architecture SYN_ARCHBEH of nd2_25266 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25265 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25265;

architecture SYN_ARCHBEH of nd2_25265 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25264 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25264;

architecture SYN_ARCHBEH of nd2_25264 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25263 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25263;

architecture SYN_ARCHBEH of nd2_25263 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25262 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25262;

architecture SYN_ARCHBEH of nd2_25262 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25261 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25261;

architecture SYN_ARCHBEH of nd2_25261 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25260 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25260;

architecture SYN_ARCHBEH of nd2_25260 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25259 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25259;

architecture SYN_ARCHBEH of nd2_25259 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25258 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25258;

architecture SYN_ARCHBEH of nd2_25258 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25257 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25257;

architecture SYN_ARCHBEH of nd2_25257 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25256 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25256;

architecture SYN_ARCHBEH of nd2_25256 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25255 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25255;

architecture SYN_ARCHBEH of nd2_25255 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25254 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25254;

architecture SYN_ARCHBEH of nd2_25254 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25253 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25253;

architecture SYN_ARCHBEH of nd2_25253 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25252 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25252;

architecture SYN_ARCHBEH of nd2_25252 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25251 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25251;

architecture SYN_ARCHBEH of nd2_25251 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25250 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25250;

architecture SYN_ARCHBEH of nd2_25250 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25249 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25249;

architecture SYN_ARCHBEH of nd2_25249 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25248 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25248;

architecture SYN_ARCHBEH of nd2_25248 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25247 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25247;

architecture SYN_ARCHBEH of nd2_25247 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25246 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25246;

architecture SYN_ARCHBEH of nd2_25246 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25245 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25245;

architecture SYN_ARCHBEH of nd2_25245 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25244 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25244;

architecture SYN_ARCHBEH of nd2_25244 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25243 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25243;

architecture SYN_ARCHBEH of nd2_25243 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25242 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25242;

architecture SYN_ARCHBEH of nd2_25242 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25241 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25241;

architecture SYN_ARCHBEH of nd2_25241 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25240 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25240;

architecture SYN_ARCHBEH of nd2_25240 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25239 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25239;

architecture SYN_ARCHBEH of nd2_25239 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25238 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25238;

architecture SYN_ARCHBEH of nd2_25238 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25237 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25237;

architecture SYN_ARCHBEH of nd2_25237 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25236 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25236;

architecture SYN_ARCHBEH of nd2_25236 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25235 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25235;

architecture SYN_ARCHBEH of nd2_25235 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25234 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25234;

architecture SYN_ARCHBEH of nd2_25234 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25233 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25233;

architecture SYN_ARCHBEH of nd2_25233 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25232 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25232;

architecture SYN_ARCHBEH of nd2_25232 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25231 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25231;

architecture SYN_ARCHBEH of nd2_25231 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25230 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25230;

architecture SYN_ARCHBEH of nd2_25230 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25229 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25229;

architecture SYN_ARCHBEH of nd2_25229 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25228 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25228;

architecture SYN_ARCHBEH of nd2_25228 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25227 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25227;

architecture SYN_ARCHBEH of nd2_25227 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25226 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25226;

architecture SYN_ARCHBEH of nd2_25226 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25225 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25225;

architecture SYN_ARCHBEH of nd2_25225 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25224 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25224;

architecture SYN_ARCHBEH of nd2_25224 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25223 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25223;

architecture SYN_ARCHBEH of nd2_25223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25222 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25222;

architecture SYN_ARCHBEH of nd2_25222 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25221 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25221;

architecture SYN_ARCHBEH of nd2_25221 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25220 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25220;

architecture SYN_ARCHBEH of nd2_25220 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25219 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25219;

architecture SYN_ARCHBEH of nd2_25219 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25218 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25218;

architecture SYN_ARCHBEH of nd2_25218 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25217 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25217;

architecture SYN_ARCHBEH of nd2_25217 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25216 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25216;

architecture SYN_ARCHBEH of nd2_25216 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25215 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25215;

architecture SYN_ARCHBEH of nd2_25215 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25214 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25214;

architecture SYN_ARCHBEH of nd2_25214 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25213 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25213;

architecture SYN_ARCHBEH of nd2_25213 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25212 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25212;

architecture SYN_ARCHBEH of nd2_25212 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25211 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25211;

architecture SYN_ARCHBEH of nd2_25211 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25210 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25210;

architecture SYN_ARCHBEH of nd2_25210 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25209 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25209;

architecture SYN_ARCHBEH of nd2_25209 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25208 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25208;

architecture SYN_ARCHBEH of nd2_25208 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25207 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25207;

architecture SYN_ARCHBEH of nd2_25207 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25206 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25206;

architecture SYN_ARCHBEH of nd2_25206 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25205 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25205;

architecture SYN_ARCHBEH of nd2_25205 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25204 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25204;

architecture SYN_ARCHBEH of nd2_25204 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25203 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25203;

architecture SYN_ARCHBEH of nd2_25203 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25202 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25202;

architecture SYN_ARCHBEH of nd2_25202 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25201 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25201;

architecture SYN_ARCHBEH of nd2_25201 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25200 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25200;

architecture SYN_ARCHBEH of nd2_25200 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25199 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25199;

architecture SYN_ARCHBEH of nd2_25199 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25198 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25198;

architecture SYN_ARCHBEH of nd2_25198 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25197 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25197;

architecture SYN_ARCHBEH of nd2_25197 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25196 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25196;

architecture SYN_ARCHBEH of nd2_25196 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25195 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25195;

architecture SYN_ARCHBEH of nd2_25195 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25194 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25194;

architecture SYN_ARCHBEH of nd2_25194 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25193 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25193;

architecture SYN_ARCHBEH of nd2_25193 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25192 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25192;

architecture SYN_ARCHBEH of nd2_25192 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25191 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25191;

architecture SYN_ARCHBEH of nd2_25191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25190 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25190;

architecture SYN_ARCHBEH of nd2_25190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25189 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25189;

architecture SYN_ARCHBEH of nd2_25189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25188 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25188;

architecture SYN_ARCHBEH of nd2_25188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25187 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25187;

architecture SYN_ARCHBEH of nd2_25187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25186 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25186;

architecture SYN_ARCHBEH of nd2_25186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25185 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25185;

architecture SYN_ARCHBEH of nd2_25185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25184 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25184;

architecture SYN_ARCHBEH of nd2_25184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25183 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25183;

architecture SYN_ARCHBEH of nd2_25183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25182 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25182;

architecture SYN_ARCHBEH of nd2_25182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25181 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25181;

architecture SYN_ARCHBEH of nd2_25181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25180 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25180;

architecture SYN_ARCHBEH of nd2_25180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25179 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25179;

architecture SYN_ARCHBEH of nd2_25179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25178 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25178;

architecture SYN_ARCHBEH of nd2_25178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25177 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25177;

architecture SYN_ARCHBEH of nd2_25177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25176 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25176;

architecture SYN_ARCHBEH of nd2_25176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25175 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25175;

architecture SYN_ARCHBEH of nd2_25175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25174 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25174;

architecture SYN_ARCHBEH of nd2_25174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25173 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25173;

architecture SYN_ARCHBEH of nd2_25173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25172 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25172;

architecture SYN_ARCHBEH of nd2_25172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25171 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25171;

architecture SYN_ARCHBEH of nd2_25171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25170 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25170;

architecture SYN_ARCHBEH of nd2_25170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25169 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25169;

architecture SYN_ARCHBEH of nd2_25169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25168 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25168;

architecture SYN_ARCHBEH of nd2_25168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25167 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25167;

architecture SYN_ARCHBEH of nd2_25167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25166 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25166;

architecture SYN_ARCHBEH of nd2_25166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25165 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25165;

architecture SYN_ARCHBEH of nd2_25165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25164 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25164;

architecture SYN_ARCHBEH of nd2_25164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25163 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25163;

architecture SYN_ARCHBEH of nd2_25163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25162 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25162;

architecture SYN_ARCHBEH of nd2_25162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25161 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25161;

architecture SYN_ARCHBEH of nd2_25161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25160 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25160;

architecture SYN_ARCHBEH of nd2_25160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25159 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25159;

architecture SYN_ARCHBEH of nd2_25159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25158 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25158;

architecture SYN_ARCHBEH of nd2_25158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25157 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25157;

architecture SYN_ARCHBEH of nd2_25157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25156 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25156;

architecture SYN_ARCHBEH of nd2_25156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25155 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25155;

architecture SYN_ARCHBEH of nd2_25155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25154 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25154;

architecture SYN_ARCHBEH of nd2_25154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25153 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25153;

architecture SYN_ARCHBEH of nd2_25153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25152 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25152;

architecture SYN_ARCHBEH of nd2_25152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25151 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25151;

architecture SYN_ARCHBEH of nd2_25151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25150 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25150;

architecture SYN_ARCHBEH of nd2_25150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25149 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25149;

architecture SYN_ARCHBEH of nd2_25149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25148 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25148;

architecture SYN_ARCHBEH of nd2_25148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25147 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25147;

architecture SYN_ARCHBEH of nd2_25147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25146 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25146;

architecture SYN_ARCHBEH of nd2_25146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25145 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25145;

architecture SYN_ARCHBEH of nd2_25145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25144 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25144;

architecture SYN_ARCHBEH of nd2_25144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25143 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25143;

architecture SYN_ARCHBEH of nd2_25143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25142 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25142;

architecture SYN_ARCHBEH of nd2_25142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25141 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25141;

architecture SYN_ARCHBEH of nd2_25141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25140 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25140;

architecture SYN_ARCHBEH of nd2_25140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25139 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25139;

architecture SYN_ARCHBEH of nd2_25139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25138 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25138;

architecture SYN_ARCHBEH of nd2_25138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25137 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25137;

architecture SYN_ARCHBEH of nd2_25137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25136 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25136;

architecture SYN_ARCHBEH of nd2_25136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25135 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25135;

architecture SYN_ARCHBEH of nd2_25135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25134 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25134;

architecture SYN_ARCHBEH of nd2_25134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25133 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25133;

architecture SYN_ARCHBEH of nd2_25133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25132 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25132;

architecture SYN_ARCHBEH of nd2_25132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25131 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25131;

architecture SYN_ARCHBEH of nd2_25131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25130 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25130;

architecture SYN_ARCHBEH of nd2_25130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25129 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25129;

architecture SYN_ARCHBEH of nd2_25129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25128 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25128;

architecture SYN_ARCHBEH of nd2_25128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25127 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25127;

architecture SYN_ARCHBEH of nd2_25127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25126 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25126;

architecture SYN_ARCHBEH of nd2_25126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25125 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25125;

architecture SYN_ARCHBEH of nd2_25125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25124 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25124;

architecture SYN_ARCHBEH of nd2_25124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25123 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25123;

architecture SYN_ARCHBEH of nd2_25123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25122 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25122;

architecture SYN_ARCHBEH of nd2_25122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25121 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25121;

architecture SYN_ARCHBEH of nd2_25121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25120 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25120;

architecture SYN_ARCHBEH of nd2_25120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25119 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25119;

architecture SYN_ARCHBEH of nd2_25119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25118 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25118;

architecture SYN_ARCHBEH of nd2_25118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25117 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25117;

architecture SYN_ARCHBEH of nd2_25117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25116 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25116;

architecture SYN_ARCHBEH of nd2_25116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25115 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25115;

architecture SYN_ARCHBEH of nd2_25115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25114 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25114;

architecture SYN_ARCHBEH of nd2_25114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25113 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25113;

architecture SYN_ARCHBEH of nd2_25113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25112 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25112;

architecture SYN_ARCHBEH of nd2_25112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25111 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25111;

architecture SYN_ARCHBEH of nd2_25111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25110 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25110;

architecture SYN_ARCHBEH of nd2_25110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25109 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25109;

architecture SYN_ARCHBEH of nd2_25109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25108 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25108;

architecture SYN_ARCHBEH of nd2_25108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25107 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25107;

architecture SYN_ARCHBEH of nd2_25107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25106 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25106;

architecture SYN_ARCHBEH of nd2_25106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25105 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25105;

architecture SYN_ARCHBEH of nd2_25105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25104 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25104;

architecture SYN_ARCHBEH of nd2_25104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25103 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25103;

architecture SYN_ARCHBEH of nd2_25103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25102 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25102;

architecture SYN_ARCHBEH of nd2_25102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25101 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25101;

architecture SYN_ARCHBEH of nd2_25101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25100 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25100;

architecture SYN_ARCHBEH of nd2_25100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25099 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25099;

architecture SYN_ARCHBEH of nd2_25099 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25098 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25098;

architecture SYN_ARCHBEH of nd2_25098 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25097 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25097;

architecture SYN_ARCHBEH of nd2_25097 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25096 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25096;

architecture SYN_ARCHBEH of nd2_25096 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25095 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25095;

architecture SYN_ARCHBEH of nd2_25095 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25094 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25094;

architecture SYN_ARCHBEH of nd2_25094 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25093 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25093;

architecture SYN_ARCHBEH of nd2_25093 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25092 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25092;

architecture SYN_ARCHBEH of nd2_25092 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25091 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25091;

architecture SYN_ARCHBEH of nd2_25091 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25090 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25090;

architecture SYN_ARCHBEH of nd2_25090 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25089 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25089;

architecture SYN_ARCHBEH of nd2_25089 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25088 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25088;

architecture SYN_ARCHBEH of nd2_25088 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25087 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25087;

architecture SYN_ARCHBEH of nd2_25087 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25086 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25086;

architecture SYN_ARCHBEH of nd2_25086 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25085 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25085;

architecture SYN_ARCHBEH of nd2_25085 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25084 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25084;

architecture SYN_ARCHBEH of nd2_25084 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25083 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25083;

architecture SYN_ARCHBEH of nd2_25083 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25082 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25082;

architecture SYN_ARCHBEH of nd2_25082 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25081 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25081;

architecture SYN_ARCHBEH of nd2_25081 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25080 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25080;

architecture SYN_ARCHBEH of nd2_25080 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25079 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25079;

architecture SYN_ARCHBEH of nd2_25079 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25078 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25078;

architecture SYN_ARCHBEH of nd2_25078 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25077 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25077;

architecture SYN_ARCHBEH of nd2_25077 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25076 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25076;

architecture SYN_ARCHBEH of nd2_25076 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25075 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25075;

architecture SYN_ARCHBEH of nd2_25075 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25074 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25074;

architecture SYN_ARCHBEH of nd2_25074 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25073 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25073;

architecture SYN_ARCHBEH of nd2_25073 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25072 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25072;

architecture SYN_ARCHBEH of nd2_25072 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25071 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25071;

architecture SYN_ARCHBEH of nd2_25071 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25070 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25070;

architecture SYN_ARCHBEH of nd2_25070 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25069 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25069;

architecture SYN_ARCHBEH of nd2_25069 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25068 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25068;

architecture SYN_ARCHBEH of nd2_25068 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25067 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25067;

architecture SYN_ARCHBEH of nd2_25067 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25066 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25066;

architecture SYN_ARCHBEH of nd2_25066 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25065 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25065;

architecture SYN_ARCHBEH of nd2_25065 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25064 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25064;

architecture SYN_ARCHBEH of nd2_25064 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25063 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25063;

architecture SYN_ARCHBEH of nd2_25063 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25062 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25062;

architecture SYN_ARCHBEH of nd2_25062 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25061 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25061;

architecture SYN_ARCHBEH of nd2_25061 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25060 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25060;

architecture SYN_ARCHBEH of nd2_25060 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25059 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25059;

architecture SYN_ARCHBEH of nd2_25059 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25058 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25058;

architecture SYN_ARCHBEH of nd2_25058 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25057 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25057;

architecture SYN_ARCHBEH of nd2_25057 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25056 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25056;

architecture SYN_ARCHBEH of nd2_25056 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25055 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25055;

architecture SYN_ARCHBEH of nd2_25055 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25054 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25054;

architecture SYN_ARCHBEH of nd2_25054 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25053 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25053;

architecture SYN_ARCHBEH of nd2_25053 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25052 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25052;

architecture SYN_ARCHBEH of nd2_25052 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25051 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25051;

architecture SYN_ARCHBEH of nd2_25051 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25050 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25050;

architecture SYN_ARCHBEH of nd2_25050 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25049 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25049;

architecture SYN_ARCHBEH of nd2_25049 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25048 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25048;

architecture SYN_ARCHBEH of nd2_25048 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25047 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25047;

architecture SYN_ARCHBEH of nd2_25047 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25046 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25046;

architecture SYN_ARCHBEH of nd2_25046 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25045 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25045;

architecture SYN_ARCHBEH of nd2_25045 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25044 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25044;

architecture SYN_ARCHBEH of nd2_25044 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25043 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25043;

architecture SYN_ARCHBEH of nd2_25043 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25042 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25042;

architecture SYN_ARCHBEH of nd2_25042 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25041 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25041;

architecture SYN_ARCHBEH of nd2_25041 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25040 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25040;

architecture SYN_ARCHBEH of nd2_25040 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25039 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25039;

architecture SYN_ARCHBEH of nd2_25039 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25038 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25038;

architecture SYN_ARCHBEH of nd2_25038 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25037 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25037;

architecture SYN_ARCHBEH of nd2_25037 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25036 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25036;

architecture SYN_ARCHBEH of nd2_25036 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25035 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25035;

architecture SYN_ARCHBEH of nd2_25035 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25034 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25034;

architecture SYN_ARCHBEH of nd2_25034 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25033 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25033;

architecture SYN_ARCHBEH of nd2_25033 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25032 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25032;

architecture SYN_ARCHBEH of nd2_25032 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25031 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25031;

architecture SYN_ARCHBEH of nd2_25031 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25030 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25030;

architecture SYN_ARCHBEH of nd2_25030 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25029 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25029;

architecture SYN_ARCHBEH of nd2_25029 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25028 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25028;

architecture SYN_ARCHBEH of nd2_25028 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25027 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25027;

architecture SYN_ARCHBEH of nd2_25027 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25026 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25026;

architecture SYN_ARCHBEH of nd2_25026 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25025 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25025;

architecture SYN_ARCHBEH of nd2_25025 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25024 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25024;

architecture SYN_ARCHBEH of nd2_25024 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25023 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25023;

architecture SYN_ARCHBEH of nd2_25023 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25022 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25022;

architecture SYN_ARCHBEH of nd2_25022 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25021 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25021;

architecture SYN_ARCHBEH of nd2_25021 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25020 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25020;

architecture SYN_ARCHBEH of nd2_25020 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25019 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25019;

architecture SYN_ARCHBEH of nd2_25019 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25018 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25018;

architecture SYN_ARCHBEH of nd2_25018 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25017 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25017;

architecture SYN_ARCHBEH of nd2_25017 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25016 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25016;

architecture SYN_ARCHBEH of nd2_25016 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25015 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25015;

architecture SYN_ARCHBEH of nd2_25015 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25014 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25014;

architecture SYN_ARCHBEH of nd2_25014 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25013 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25013;

architecture SYN_ARCHBEH of nd2_25013 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25012 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25012;

architecture SYN_ARCHBEH of nd2_25012 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25011 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25011;

architecture SYN_ARCHBEH of nd2_25011 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25010 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25010;

architecture SYN_ARCHBEH of nd2_25010 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25009 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25009;

architecture SYN_ARCHBEH of nd2_25009 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25008 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25008;

architecture SYN_ARCHBEH of nd2_25008 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25007 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25007;

architecture SYN_ARCHBEH of nd2_25007 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25006 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25006;

architecture SYN_ARCHBEH of nd2_25006 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25005 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25005;

architecture SYN_ARCHBEH of nd2_25005 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25004 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25004;

architecture SYN_ARCHBEH of nd2_25004 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25003 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25003;

architecture SYN_ARCHBEH of nd2_25003 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25002 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25002;

architecture SYN_ARCHBEH of nd2_25002 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25001 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25001;

architecture SYN_ARCHBEH of nd2_25001 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_25000 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_25000;

architecture SYN_ARCHBEH of nd2_25000 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24999 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24999;

architecture SYN_ARCHBEH of nd2_24999 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24998 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24998;

architecture SYN_ARCHBEH of nd2_24998 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24997 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24997;

architecture SYN_ARCHBEH of nd2_24997 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24996 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24996;

architecture SYN_ARCHBEH of nd2_24996 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24995 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24995;

architecture SYN_ARCHBEH of nd2_24995 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24994 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24994;

architecture SYN_ARCHBEH of nd2_24994 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24993 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24993;

architecture SYN_ARCHBEH of nd2_24993 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24992 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24992;

architecture SYN_ARCHBEH of nd2_24992 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24991 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24991;

architecture SYN_ARCHBEH of nd2_24991 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24990 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24990;

architecture SYN_ARCHBEH of nd2_24990 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24989 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24989;

architecture SYN_ARCHBEH of nd2_24989 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24988 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24988;

architecture SYN_ARCHBEH of nd2_24988 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24987 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24987;

architecture SYN_ARCHBEH of nd2_24987 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24986 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24986;

architecture SYN_ARCHBEH of nd2_24986 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24985 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24985;

architecture SYN_ARCHBEH of nd2_24985 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24984 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24984;

architecture SYN_ARCHBEH of nd2_24984 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24983 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24983;

architecture SYN_ARCHBEH of nd2_24983 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24982 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24982;

architecture SYN_ARCHBEH of nd2_24982 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24981 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24981;

architecture SYN_ARCHBEH of nd2_24981 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24980 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24980;

architecture SYN_ARCHBEH of nd2_24980 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24979 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24979;

architecture SYN_ARCHBEH of nd2_24979 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24978 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24978;

architecture SYN_ARCHBEH of nd2_24978 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24977 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24977;

architecture SYN_ARCHBEH of nd2_24977 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24976 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24976;

architecture SYN_ARCHBEH of nd2_24976 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24975 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24975;

architecture SYN_ARCHBEH of nd2_24975 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24974 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24974;

architecture SYN_ARCHBEH of nd2_24974 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24973 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24973;

architecture SYN_ARCHBEH of nd2_24973 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24972 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24972;

architecture SYN_ARCHBEH of nd2_24972 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24971 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24971;

architecture SYN_ARCHBEH of nd2_24971 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24970 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24970;

architecture SYN_ARCHBEH of nd2_24970 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24969 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24969;

architecture SYN_ARCHBEH of nd2_24969 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24968 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24968;

architecture SYN_ARCHBEH of nd2_24968 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24967 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24967;

architecture SYN_ARCHBEH of nd2_24967 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24966 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24966;

architecture SYN_ARCHBEH of nd2_24966 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24965 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24965;

architecture SYN_ARCHBEH of nd2_24965 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24964 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24964;

architecture SYN_ARCHBEH of nd2_24964 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24963 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24963;

architecture SYN_ARCHBEH of nd2_24963 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24962 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24962;

architecture SYN_ARCHBEH of nd2_24962 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24961 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24961;

architecture SYN_ARCHBEH of nd2_24961 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24960 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24960;

architecture SYN_ARCHBEH of nd2_24960 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24959 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24959;

architecture SYN_ARCHBEH of nd2_24959 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24958 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24958;

architecture SYN_ARCHBEH of nd2_24958 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24957 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24957;

architecture SYN_ARCHBEH of nd2_24957 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24956 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24956;

architecture SYN_ARCHBEH of nd2_24956 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24955 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24955;

architecture SYN_ARCHBEH of nd2_24955 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24954 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24954;

architecture SYN_ARCHBEH of nd2_24954 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24953 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24953;

architecture SYN_ARCHBEH of nd2_24953 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24952 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24952;

architecture SYN_ARCHBEH of nd2_24952 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24951 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24951;

architecture SYN_ARCHBEH of nd2_24951 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24950 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24950;

architecture SYN_ARCHBEH of nd2_24950 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24949 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24949;

architecture SYN_ARCHBEH of nd2_24949 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24948 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24948;

architecture SYN_ARCHBEH of nd2_24948 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24947 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24947;

architecture SYN_ARCHBEH of nd2_24947 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24946 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24946;

architecture SYN_ARCHBEH of nd2_24946 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24945 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24945;

architecture SYN_ARCHBEH of nd2_24945 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24944 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24944;

architecture SYN_ARCHBEH of nd2_24944 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24943 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24943;

architecture SYN_ARCHBEH of nd2_24943 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24942 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24942;

architecture SYN_ARCHBEH of nd2_24942 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24941 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24941;

architecture SYN_ARCHBEH of nd2_24941 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24940 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24940;

architecture SYN_ARCHBEH of nd2_24940 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24939 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24939;

architecture SYN_ARCHBEH of nd2_24939 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24938 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24938;

architecture SYN_ARCHBEH of nd2_24938 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24937 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24937;

architecture SYN_ARCHBEH of nd2_24937 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24936 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24936;

architecture SYN_ARCHBEH of nd2_24936 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24935 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24935;

architecture SYN_ARCHBEH of nd2_24935 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24934 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24934;

architecture SYN_ARCHBEH of nd2_24934 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24933 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24933;

architecture SYN_ARCHBEH of nd2_24933 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24932 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24932;

architecture SYN_ARCHBEH of nd2_24932 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24931 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24931;

architecture SYN_ARCHBEH of nd2_24931 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24930 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24930;

architecture SYN_ARCHBEH of nd2_24930 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24929 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24929;

architecture SYN_ARCHBEH of nd2_24929 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24928 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24928;

architecture SYN_ARCHBEH of nd2_24928 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24927 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24927;

architecture SYN_ARCHBEH of nd2_24927 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24926 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24926;

architecture SYN_ARCHBEH of nd2_24926 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24925 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24925;

architecture SYN_ARCHBEH of nd2_24925 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24924 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24924;

architecture SYN_ARCHBEH of nd2_24924 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24923 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24923;

architecture SYN_ARCHBEH of nd2_24923 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24922 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24922;

architecture SYN_ARCHBEH of nd2_24922 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24921 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24921;

architecture SYN_ARCHBEH of nd2_24921 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24920 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24920;

architecture SYN_ARCHBEH of nd2_24920 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24919 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24919;

architecture SYN_ARCHBEH of nd2_24919 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24918 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24918;

architecture SYN_ARCHBEH of nd2_24918 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24917 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24917;

architecture SYN_ARCHBEH of nd2_24917 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24916 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24916;

architecture SYN_ARCHBEH of nd2_24916 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24915 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24915;

architecture SYN_ARCHBEH of nd2_24915 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24914 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24914;

architecture SYN_ARCHBEH of nd2_24914 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24913 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24913;

architecture SYN_ARCHBEH of nd2_24913 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24912 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24912;

architecture SYN_ARCHBEH of nd2_24912 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24911 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24911;

architecture SYN_ARCHBEH of nd2_24911 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24910 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24910;

architecture SYN_ARCHBEH of nd2_24910 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24909 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24909;

architecture SYN_ARCHBEH of nd2_24909 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24908 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24908;

architecture SYN_ARCHBEH of nd2_24908 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24907 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24907;

architecture SYN_ARCHBEH of nd2_24907 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24906 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24906;

architecture SYN_ARCHBEH of nd2_24906 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24905 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24905;

architecture SYN_ARCHBEH of nd2_24905 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24904 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24904;

architecture SYN_ARCHBEH of nd2_24904 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24903 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24903;

architecture SYN_ARCHBEH of nd2_24903 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24902 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24902;

architecture SYN_ARCHBEH of nd2_24902 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24901 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24901;

architecture SYN_ARCHBEH of nd2_24901 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24900 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24900;

architecture SYN_ARCHBEH of nd2_24900 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24899 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24899;

architecture SYN_ARCHBEH of nd2_24899 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24898 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24898;

architecture SYN_ARCHBEH of nd2_24898 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24897 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24897;

architecture SYN_ARCHBEH of nd2_24897 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24896 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24896;

architecture SYN_ARCHBEH of nd2_24896 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24895 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24895;

architecture SYN_ARCHBEH of nd2_24895 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24894 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24894;

architecture SYN_ARCHBEH of nd2_24894 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24893 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24893;

architecture SYN_ARCHBEH of nd2_24893 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24892 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24892;

architecture SYN_ARCHBEH of nd2_24892 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24891 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24891;

architecture SYN_ARCHBEH of nd2_24891 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24890 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24890;

architecture SYN_ARCHBEH of nd2_24890 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24889 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24889;

architecture SYN_ARCHBEH of nd2_24889 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24888 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24888;

architecture SYN_ARCHBEH of nd2_24888 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24887 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24887;

architecture SYN_ARCHBEH of nd2_24887 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24886 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24886;

architecture SYN_ARCHBEH of nd2_24886 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24885 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24885;

architecture SYN_ARCHBEH of nd2_24885 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24884 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24884;

architecture SYN_ARCHBEH of nd2_24884 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24883 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24883;

architecture SYN_ARCHBEH of nd2_24883 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24882 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24882;

architecture SYN_ARCHBEH of nd2_24882 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24881 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24881;

architecture SYN_ARCHBEH of nd2_24881 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24880 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24880;

architecture SYN_ARCHBEH of nd2_24880 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24879 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24879;

architecture SYN_ARCHBEH of nd2_24879 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24878 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24878;

architecture SYN_ARCHBEH of nd2_24878 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24877 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24877;

architecture SYN_ARCHBEH of nd2_24877 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24876 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24876;

architecture SYN_ARCHBEH of nd2_24876 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24875 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24875;

architecture SYN_ARCHBEH of nd2_24875 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24874 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24874;

architecture SYN_ARCHBEH of nd2_24874 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24873 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24873;

architecture SYN_ARCHBEH of nd2_24873 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24872 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24872;

architecture SYN_ARCHBEH of nd2_24872 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24871 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24871;

architecture SYN_ARCHBEH of nd2_24871 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24870 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24870;

architecture SYN_ARCHBEH of nd2_24870 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24869 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24869;

architecture SYN_ARCHBEH of nd2_24869 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24868 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24868;

architecture SYN_ARCHBEH of nd2_24868 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24867 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24867;

architecture SYN_ARCHBEH of nd2_24867 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24866 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24866;

architecture SYN_ARCHBEH of nd2_24866 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24865 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24865;

architecture SYN_ARCHBEH of nd2_24865 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24864 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24864;

architecture SYN_ARCHBEH of nd2_24864 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24863 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24863;

architecture SYN_ARCHBEH of nd2_24863 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24862 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24862;

architecture SYN_ARCHBEH of nd2_24862 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24861 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24861;

architecture SYN_ARCHBEH of nd2_24861 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24860 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24860;

architecture SYN_ARCHBEH of nd2_24860 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24859 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24859;

architecture SYN_ARCHBEH of nd2_24859 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24858 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24858;

architecture SYN_ARCHBEH of nd2_24858 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24857 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24857;

architecture SYN_ARCHBEH of nd2_24857 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24856 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24856;

architecture SYN_ARCHBEH of nd2_24856 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24855 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24855;

architecture SYN_ARCHBEH of nd2_24855 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24854 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24854;

architecture SYN_ARCHBEH of nd2_24854 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24853 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24853;

architecture SYN_ARCHBEH of nd2_24853 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24852 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24852;

architecture SYN_ARCHBEH of nd2_24852 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24851 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24851;

architecture SYN_ARCHBEH of nd2_24851 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24850 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24850;

architecture SYN_ARCHBEH of nd2_24850 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24849 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24849;

architecture SYN_ARCHBEH of nd2_24849 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24848 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24848;

architecture SYN_ARCHBEH of nd2_24848 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24847 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24847;

architecture SYN_ARCHBEH of nd2_24847 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24846 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24846;

architecture SYN_ARCHBEH of nd2_24846 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24845 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24845;

architecture SYN_ARCHBEH of nd2_24845 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24844 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24844;

architecture SYN_ARCHBEH of nd2_24844 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24843 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24843;

architecture SYN_ARCHBEH of nd2_24843 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24842 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24842;

architecture SYN_ARCHBEH of nd2_24842 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24841 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24841;

architecture SYN_ARCHBEH of nd2_24841 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24840 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24840;

architecture SYN_ARCHBEH of nd2_24840 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24839 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24839;

architecture SYN_ARCHBEH of nd2_24839 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24838 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24838;

architecture SYN_ARCHBEH of nd2_24838 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24837 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24837;

architecture SYN_ARCHBEH of nd2_24837 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24836 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24836;

architecture SYN_ARCHBEH of nd2_24836 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24835 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24835;

architecture SYN_ARCHBEH of nd2_24835 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24834 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24834;

architecture SYN_ARCHBEH of nd2_24834 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24833 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24833;

architecture SYN_ARCHBEH of nd2_24833 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24832 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24832;

architecture SYN_ARCHBEH of nd2_24832 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24831 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24831;

architecture SYN_ARCHBEH of nd2_24831 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24830 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24830;

architecture SYN_ARCHBEH of nd2_24830 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24829 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24829;

architecture SYN_ARCHBEH of nd2_24829 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24828 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24828;

architecture SYN_ARCHBEH of nd2_24828 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24827 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24827;

architecture SYN_ARCHBEH of nd2_24827 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24826 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24826;

architecture SYN_ARCHBEH of nd2_24826 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24825 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24825;

architecture SYN_ARCHBEH of nd2_24825 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24824 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24824;

architecture SYN_ARCHBEH of nd2_24824 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24823 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24823;

architecture SYN_ARCHBEH of nd2_24823 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24822 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24822;

architecture SYN_ARCHBEH of nd2_24822 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24821 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24821;

architecture SYN_ARCHBEH of nd2_24821 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24820 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24820;

architecture SYN_ARCHBEH of nd2_24820 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24819 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24819;

architecture SYN_ARCHBEH of nd2_24819 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24818 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24818;

architecture SYN_ARCHBEH of nd2_24818 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24817 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24817;

architecture SYN_ARCHBEH of nd2_24817 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24816 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24816;

architecture SYN_ARCHBEH of nd2_24816 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24815 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24815;

architecture SYN_ARCHBEH of nd2_24815 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24814 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24814;

architecture SYN_ARCHBEH of nd2_24814 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24813 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24813;

architecture SYN_ARCHBEH of nd2_24813 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24812 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24812;

architecture SYN_ARCHBEH of nd2_24812 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24811 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24811;

architecture SYN_ARCHBEH of nd2_24811 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24810 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24810;

architecture SYN_ARCHBEH of nd2_24810 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24809 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24809;

architecture SYN_ARCHBEH of nd2_24809 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24808 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24808;

architecture SYN_ARCHBEH of nd2_24808 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24807 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24807;

architecture SYN_ARCHBEH of nd2_24807 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24806 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24806;

architecture SYN_ARCHBEH of nd2_24806 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24805 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24805;

architecture SYN_ARCHBEH of nd2_24805 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24804 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24804;

architecture SYN_ARCHBEH of nd2_24804 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24803 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24803;

architecture SYN_ARCHBEH of nd2_24803 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24802 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24802;

architecture SYN_ARCHBEH of nd2_24802 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24801 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24801;

architecture SYN_ARCHBEH of nd2_24801 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24800 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24800;

architecture SYN_ARCHBEH of nd2_24800 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24799 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24799;

architecture SYN_ARCHBEH of nd2_24799 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24798 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24798;

architecture SYN_ARCHBEH of nd2_24798 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24797 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24797;

architecture SYN_ARCHBEH of nd2_24797 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24796 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24796;

architecture SYN_ARCHBEH of nd2_24796 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24795 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24795;

architecture SYN_ARCHBEH of nd2_24795 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24794 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24794;

architecture SYN_ARCHBEH of nd2_24794 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24793 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24793;

architecture SYN_ARCHBEH of nd2_24793 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24792 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24792;

architecture SYN_ARCHBEH of nd2_24792 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24791 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24791;

architecture SYN_ARCHBEH of nd2_24791 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24790 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24790;

architecture SYN_ARCHBEH of nd2_24790 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24789 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24789;

architecture SYN_ARCHBEH of nd2_24789 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24788 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24788;

architecture SYN_ARCHBEH of nd2_24788 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24787 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24787;

architecture SYN_ARCHBEH of nd2_24787 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24786 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24786;

architecture SYN_ARCHBEH of nd2_24786 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24785 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24785;

architecture SYN_ARCHBEH of nd2_24785 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24784 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24784;

architecture SYN_ARCHBEH of nd2_24784 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24783 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24783;

architecture SYN_ARCHBEH of nd2_24783 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24782 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24782;

architecture SYN_ARCHBEH of nd2_24782 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24781 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24781;

architecture SYN_ARCHBEH of nd2_24781 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24780 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24780;

architecture SYN_ARCHBEH of nd2_24780 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24779 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24779;

architecture SYN_ARCHBEH of nd2_24779 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24778 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24778;

architecture SYN_ARCHBEH of nd2_24778 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24777 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24777;

architecture SYN_ARCHBEH of nd2_24777 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24776 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24776;

architecture SYN_ARCHBEH of nd2_24776 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24775 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24775;

architecture SYN_ARCHBEH of nd2_24775 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24774 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24774;

architecture SYN_ARCHBEH of nd2_24774 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24773 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24773;

architecture SYN_ARCHBEH of nd2_24773 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24772 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24772;

architecture SYN_ARCHBEH of nd2_24772 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24771 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24771;

architecture SYN_ARCHBEH of nd2_24771 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24770 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24770;

architecture SYN_ARCHBEH of nd2_24770 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24769 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24769;

architecture SYN_ARCHBEH of nd2_24769 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24768 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24768;

architecture SYN_ARCHBEH of nd2_24768 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24767 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24767;

architecture SYN_ARCHBEH of nd2_24767 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24766 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24766;

architecture SYN_ARCHBEH of nd2_24766 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24765 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24765;

architecture SYN_ARCHBEH of nd2_24765 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24764 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24764;

architecture SYN_ARCHBEH of nd2_24764 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24763 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24763;

architecture SYN_ARCHBEH of nd2_24763 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24762 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24762;

architecture SYN_ARCHBEH of nd2_24762 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24761 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24761;

architecture SYN_ARCHBEH of nd2_24761 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24760 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24760;

architecture SYN_ARCHBEH of nd2_24760 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24759 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24759;

architecture SYN_ARCHBEH of nd2_24759 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24758 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24758;

architecture SYN_ARCHBEH of nd2_24758 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24757 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24757;

architecture SYN_ARCHBEH of nd2_24757 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24756 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24756;

architecture SYN_ARCHBEH of nd2_24756 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24755 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24755;

architecture SYN_ARCHBEH of nd2_24755 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24754 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24754;

architecture SYN_ARCHBEH of nd2_24754 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24753 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24753;

architecture SYN_ARCHBEH of nd2_24753 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24752 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24752;

architecture SYN_ARCHBEH of nd2_24752 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24751 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24751;

architecture SYN_ARCHBEH of nd2_24751 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24750 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24750;

architecture SYN_ARCHBEH of nd2_24750 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24749 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24749;

architecture SYN_ARCHBEH of nd2_24749 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24748 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24748;

architecture SYN_ARCHBEH of nd2_24748 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24747 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24747;

architecture SYN_ARCHBEH of nd2_24747 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24746 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24746;

architecture SYN_ARCHBEH of nd2_24746 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24745 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24745;

architecture SYN_ARCHBEH of nd2_24745 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24744 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24744;

architecture SYN_ARCHBEH of nd2_24744 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24743 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24743;

architecture SYN_ARCHBEH of nd2_24743 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24742 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24742;

architecture SYN_ARCHBEH of nd2_24742 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24741 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24741;

architecture SYN_ARCHBEH of nd2_24741 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24740 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24740;

architecture SYN_ARCHBEH of nd2_24740 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24739 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24739;

architecture SYN_ARCHBEH of nd2_24739 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24738 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24738;

architecture SYN_ARCHBEH of nd2_24738 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24737 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24737;

architecture SYN_ARCHBEH of nd2_24737 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24736 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24736;

architecture SYN_ARCHBEH of nd2_24736 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24735 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24735;

architecture SYN_ARCHBEH of nd2_24735 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24734 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24734;

architecture SYN_ARCHBEH of nd2_24734 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24733 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24733;

architecture SYN_ARCHBEH of nd2_24733 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24732 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24732;

architecture SYN_ARCHBEH of nd2_24732 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24731 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24731;

architecture SYN_ARCHBEH of nd2_24731 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24730 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24730;

architecture SYN_ARCHBEH of nd2_24730 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24729 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24729;

architecture SYN_ARCHBEH of nd2_24729 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24728 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24728;

architecture SYN_ARCHBEH of nd2_24728 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24727 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24727;

architecture SYN_ARCHBEH of nd2_24727 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24726 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24726;

architecture SYN_ARCHBEH of nd2_24726 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24725 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24725;

architecture SYN_ARCHBEH of nd2_24725 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24724 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24724;

architecture SYN_ARCHBEH of nd2_24724 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24723 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24723;

architecture SYN_ARCHBEH of nd2_24723 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24722 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24722;

architecture SYN_ARCHBEH of nd2_24722 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24721 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24721;

architecture SYN_ARCHBEH of nd2_24721 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24720 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24720;

architecture SYN_ARCHBEH of nd2_24720 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24719 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24719;

architecture SYN_ARCHBEH of nd2_24719 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24718 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24718;

architecture SYN_ARCHBEH of nd2_24718 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24717 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24717;

architecture SYN_ARCHBEH of nd2_24717 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24716 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24716;

architecture SYN_ARCHBEH of nd2_24716 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24715 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24715;

architecture SYN_ARCHBEH of nd2_24715 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24714 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24714;

architecture SYN_ARCHBEH of nd2_24714 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24713 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24713;

architecture SYN_ARCHBEH of nd2_24713 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24712 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24712;

architecture SYN_ARCHBEH of nd2_24712 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24711 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24711;

architecture SYN_ARCHBEH of nd2_24711 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24710 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24710;

architecture SYN_ARCHBEH of nd2_24710 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24709 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24709;

architecture SYN_ARCHBEH of nd2_24709 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24708 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24708;

architecture SYN_ARCHBEH of nd2_24708 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24707 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24707;

architecture SYN_ARCHBEH of nd2_24707 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24706 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24706;

architecture SYN_ARCHBEH of nd2_24706 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24705 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24705;

architecture SYN_ARCHBEH of nd2_24705 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24704 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24704;

architecture SYN_ARCHBEH of nd2_24704 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24703 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24703;

architecture SYN_ARCHBEH of nd2_24703 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24702 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24702;

architecture SYN_ARCHBEH of nd2_24702 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24701 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24701;

architecture SYN_ARCHBEH of nd2_24701 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24700 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24700;

architecture SYN_ARCHBEH of nd2_24700 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24699 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24699;

architecture SYN_ARCHBEH of nd2_24699 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24698 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24698;

architecture SYN_ARCHBEH of nd2_24698 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24697 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24697;

architecture SYN_ARCHBEH of nd2_24697 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24696 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24696;

architecture SYN_ARCHBEH of nd2_24696 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24695 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24695;

architecture SYN_ARCHBEH of nd2_24695 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24694 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24694;

architecture SYN_ARCHBEH of nd2_24694 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24693 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24693;

architecture SYN_ARCHBEH of nd2_24693 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24692 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24692;

architecture SYN_ARCHBEH of nd2_24692 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24691 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24691;

architecture SYN_ARCHBEH of nd2_24691 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24690 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24690;

architecture SYN_ARCHBEH of nd2_24690 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24689 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24689;

architecture SYN_ARCHBEH of nd2_24689 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24688 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24688;

architecture SYN_ARCHBEH of nd2_24688 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24687 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24687;

architecture SYN_ARCHBEH of nd2_24687 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24686 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24686;

architecture SYN_ARCHBEH of nd2_24686 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24685 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24685;

architecture SYN_ARCHBEH of nd2_24685 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24684 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24684;

architecture SYN_ARCHBEH of nd2_24684 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24683 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24683;

architecture SYN_ARCHBEH of nd2_24683 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24682 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24682;

architecture SYN_ARCHBEH of nd2_24682 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24681 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24681;

architecture SYN_ARCHBEH of nd2_24681 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24680 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24680;

architecture SYN_ARCHBEH of nd2_24680 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24679 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24679;

architecture SYN_ARCHBEH of nd2_24679 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24678 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24678;

architecture SYN_ARCHBEH of nd2_24678 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24677 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24677;

architecture SYN_ARCHBEH of nd2_24677 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24676 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24676;

architecture SYN_ARCHBEH of nd2_24676 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24675 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24675;

architecture SYN_ARCHBEH of nd2_24675 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24674 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24674;

architecture SYN_ARCHBEH of nd2_24674 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24673 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24673;

architecture SYN_ARCHBEH of nd2_24673 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24672 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24672;

architecture SYN_ARCHBEH of nd2_24672 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24671 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24671;

architecture SYN_ARCHBEH of nd2_24671 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24670 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24670;

architecture SYN_ARCHBEH of nd2_24670 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24669 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24669;

architecture SYN_ARCHBEH of nd2_24669 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24668 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24668;

architecture SYN_ARCHBEH of nd2_24668 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24667 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24667;

architecture SYN_ARCHBEH of nd2_24667 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24666 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24666;

architecture SYN_ARCHBEH of nd2_24666 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24665 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24665;

architecture SYN_ARCHBEH of nd2_24665 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24664 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24664;

architecture SYN_ARCHBEH of nd2_24664 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24663 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24663;

architecture SYN_ARCHBEH of nd2_24663 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24662 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24662;

architecture SYN_ARCHBEH of nd2_24662 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24661 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24661;

architecture SYN_ARCHBEH of nd2_24661 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24660 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24660;

architecture SYN_ARCHBEH of nd2_24660 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24659 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24659;

architecture SYN_ARCHBEH of nd2_24659 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24658 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24658;

architecture SYN_ARCHBEH of nd2_24658 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24657 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24657;

architecture SYN_ARCHBEH of nd2_24657 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24656 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24656;

architecture SYN_ARCHBEH of nd2_24656 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24655 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24655;

architecture SYN_ARCHBEH of nd2_24655 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24654 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24654;

architecture SYN_ARCHBEH of nd2_24654 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24653 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24653;

architecture SYN_ARCHBEH of nd2_24653 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24652 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24652;

architecture SYN_ARCHBEH of nd2_24652 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24651 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24651;

architecture SYN_ARCHBEH of nd2_24651 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24650 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24650;

architecture SYN_ARCHBEH of nd2_24650 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24649 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24649;

architecture SYN_ARCHBEH of nd2_24649 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24648 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24648;

architecture SYN_ARCHBEH of nd2_24648 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24647 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24647;

architecture SYN_ARCHBEH of nd2_24647 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24646 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24646;

architecture SYN_ARCHBEH of nd2_24646 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24645 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24645;

architecture SYN_ARCHBEH of nd2_24645 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24644 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24644;

architecture SYN_ARCHBEH of nd2_24644 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24643 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24643;

architecture SYN_ARCHBEH of nd2_24643 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24642 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24642;

architecture SYN_ARCHBEH of nd2_24642 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24641 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24641;

architecture SYN_ARCHBEH of nd2_24641 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24640 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24640;

architecture SYN_ARCHBEH of nd2_24640 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24639 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24639;

architecture SYN_ARCHBEH of nd2_24639 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24638 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24638;

architecture SYN_ARCHBEH of nd2_24638 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24637 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24637;

architecture SYN_ARCHBEH of nd2_24637 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24636 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24636;

architecture SYN_ARCHBEH of nd2_24636 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24635 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24635;

architecture SYN_ARCHBEH of nd2_24635 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24634 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24634;

architecture SYN_ARCHBEH of nd2_24634 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24633 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24633;

architecture SYN_ARCHBEH of nd2_24633 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24632 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24632;

architecture SYN_ARCHBEH of nd2_24632 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24631 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24631;

architecture SYN_ARCHBEH of nd2_24631 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24630 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24630;

architecture SYN_ARCHBEH of nd2_24630 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24629 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24629;

architecture SYN_ARCHBEH of nd2_24629 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24628 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24628;

architecture SYN_ARCHBEH of nd2_24628 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24627 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24627;

architecture SYN_ARCHBEH of nd2_24627 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24626 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24626;

architecture SYN_ARCHBEH of nd2_24626 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24625 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24625;

architecture SYN_ARCHBEH of nd2_24625 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24624 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24624;

architecture SYN_ARCHBEH of nd2_24624 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24623 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24623;

architecture SYN_ARCHBEH of nd2_24623 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24622 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24622;

architecture SYN_ARCHBEH of nd2_24622 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24621 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24621;

architecture SYN_ARCHBEH of nd2_24621 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24620 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24620;

architecture SYN_ARCHBEH of nd2_24620 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24619 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24619;

architecture SYN_ARCHBEH of nd2_24619 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24618 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24618;

architecture SYN_ARCHBEH of nd2_24618 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24617 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24617;

architecture SYN_ARCHBEH of nd2_24617 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24616 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24616;

architecture SYN_ARCHBEH of nd2_24616 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24615 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24615;

architecture SYN_ARCHBEH of nd2_24615 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24614 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24614;

architecture SYN_ARCHBEH of nd2_24614 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24613 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24613;

architecture SYN_ARCHBEH of nd2_24613 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24612 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24612;

architecture SYN_ARCHBEH of nd2_24612 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24611 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24611;

architecture SYN_ARCHBEH of nd2_24611 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24610 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24610;

architecture SYN_ARCHBEH of nd2_24610 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24609 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24609;

architecture SYN_ARCHBEH of nd2_24609 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24608 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24608;

architecture SYN_ARCHBEH of nd2_24608 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24607 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24607;

architecture SYN_ARCHBEH of nd2_24607 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24606 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24606;

architecture SYN_ARCHBEH of nd2_24606 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24605 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24605;

architecture SYN_ARCHBEH of nd2_24605 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24604 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24604;

architecture SYN_ARCHBEH of nd2_24604 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24603 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24603;

architecture SYN_ARCHBEH of nd2_24603 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24602 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24602;

architecture SYN_ARCHBEH of nd2_24602 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24601 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24601;

architecture SYN_ARCHBEH of nd2_24601 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24600 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24600;

architecture SYN_ARCHBEH of nd2_24600 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24599 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24599;

architecture SYN_ARCHBEH of nd2_24599 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24598 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24598;

architecture SYN_ARCHBEH of nd2_24598 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24597 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24597;

architecture SYN_ARCHBEH of nd2_24597 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24596 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24596;

architecture SYN_ARCHBEH of nd2_24596 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24595 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24595;

architecture SYN_ARCHBEH of nd2_24595 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24594 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24594;

architecture SYN_ARCHBEH of nd2_24594 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24593 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24593;

architecture SYN_ARCHBEH of nd2_24593 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24592 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24592;

architecture SYN_ARCHBEH of nd2_24592 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24591 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24591;

architecture SYN_ARCHBEH of nd2_24591 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24590 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24590;

architecture SYN_ARCHBEH of nd2_24590 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24589 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24589;

architecture SYN_ARCHBEH of nd2_24589 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24588 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24588;

architecture SYN_ARCHBEH of nd2_24588 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24587 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24587;

architecture SYN_ARCHBEH of nd2_24587 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24586 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24586;

architecture SYN_ARCHBEH of nd2_24586 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24585 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24585;

architecture SYN_ARCHBEH of nd2_24585 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24584 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24584;

architecture SYN_ARCHBEH of nd2_24584 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24583 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24583;

architecture SYN_ARCHBEH of nd2_24583 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24582 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24582;

architecture SYN_ARCHBEH of nd2_24582 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24581 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24581;

architecture SYN_ARCHBEH of nd2_24581 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24580 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24580;

architecture SYN_ARCHBEH of nd2_24580 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24579 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24579;

architecture SYN_ARCHBEH of nd2_24579 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24578 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24578;

architecture SYN_ARCHBEH of nd2_24578 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24577 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24577;

architecture SYN_ARCHBEH of nd2_24577 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24576 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24576;

architecture SYN_ARCHBEH of nd2_24576 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24575 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24575;

architecture SYN_ARCHBEH of nd2_24575 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24574 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24574;

architecture SYN_ARCHBEH of nd2_24574 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24573 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24573;

architecture SYN_ARCHBEH of nd2_24573 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24572 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24572;

architecture SYN_ARCHBEH of nd2_24572 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24571 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24571;

architecture SYN_ARCHBEH of nd2_24571 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24570 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24570;

architecture SYN_ARCHBEH of nd2_24570 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24569 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24569;

architecture SYN_ARCHBEH of nd2_24569 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24568 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24568;

architecture SYN_ARCHBEH of nd2_24568 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24567 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24567;

architecture SYN_ARCHBEH of nd2_24567 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24566 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24566;

architecture SYN_ARCHBEH of nd2_24566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24565 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24565;

architecture SYN_ARCHBEH of nd2_24565 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24564 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24564;

architecture SYN_ARCHBEH of nd2_24564 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24563 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24563;

architecture SYN_ARCHBEH of nd2_24563 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24562 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24562;

architecture SYN_ARCHBEH of nd2_24562 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24561 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24561;

architecture SYN_ARCHBEH of nd2_24561 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24560 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24560;

architecture SYN_ARCHBEH of nd2_24560 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24559 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24559;

architecture SYN_ARCHBEH of nd2_24559 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24558 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24558;

architecture SYN_ARCHBEH of nd2_24558 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24557 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24557;

architecture SYN_ARCHBEH of nd2_24557 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24556 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24556;

architecture SYN_ARCHBEH of nd2_24556 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24555 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24555;

architecture SYN_ARCHBEH of nd2_24555 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24554 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24554;

architecture SYN_ARCHBEH of nd2_24554 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24553 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24553;

architecture SYN_ARCHBEH of nd2_24553 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24552 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24552;

architecture SYN_ARCHBEH of nd2_24552 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24551 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24551;

architecture SYN_ARCHBEH of nd2_24551 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24550 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24550;

architecture SYN_ARCHBEH of nd2_24550 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24549 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24549;

architecture SYN_ARCHBEH of nd2_24549 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24548 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24548;

architecture SYN_ARCHBEH of nd2_24548 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24547 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24547;

architecture SYN_ARCHBEH of nd2_24547 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24546 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24546;

architecture SYN_ARCHBEH of nd2_24546 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24545 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24545;

architecture SYN_ARCHBEH of nd2_24545 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24544 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24544;

architecture SYN_ARCHBEH of nd2_24544 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24543 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24543;

architecture SYN_ARCHBEH of nd2_24543 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24542 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24542;

architecture SYN_ARCHBEH of nd2_24542 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24541 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24541;

architecture SYN_ARCHBEH of nd2_24541 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24540 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24540;

architecture SYN_ARCHBEH of nd2_24540 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24539 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24539;

architecture SYN_ARCHBEH of nd2_24539 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24538 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24538;

architecture SYN_ARCHBEH of nd2_24538 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24537 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24537;

architecture SYN_ARCHBEH of nd2_24537 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24536 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24536;

architecture SYN_ARCHBEH of nd2_24536 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24535 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24535;

architecture SYN_ARCHBEH of nd2_24535 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24534 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24534;

architecture SYN_ARCHBEH of nd2_24534 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24533 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24533;

architecture SYN_ARCHBEH of nd2_24533 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24532 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24532;

architecture SYN_ARCHBEH of nd2_24532 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24531 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24531;

architecture SYN_ARCHBEH of nd2_24531 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24530 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24530;

architecture SYN_ARCHBEH of nd2_24530 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24529 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24529;

architecture SYN_ARCHBEH of nd2_24529 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24528 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24528;

architecture SYN_ARCHBEH of nd2_24528 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24527 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24527;

architecture SYN_ARCHBEH of nd2_24527 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24526 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24526;

architecture SYN_ARCHBEH of nd2_24526 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24525 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24525;

architecture SYN_ARCHBEH of nd2_24525 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24524 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24524;

architecture SYN_ARCHBEH of nd2_24524 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24523 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24523;

architecture SYN_ARCHBEH of nd2_24523 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24522 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24522;

architecture SYN_ARCHBEH of nd2_24522 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24521 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24521;

architecture SYN_ARCHBEH of nd2_24521 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24520 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24520;

architecture SYN_ARCHBEH of nd2_24520 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24519 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24519;

architecture SYN_ARCHBEH of nd2_24519 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24518 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24518;

architecture SYN_ARCHBEH of nd2_24518 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24517 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24517;

architecture SYN_ARCHBEH of nd2_24517 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24516 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24516;

architecture SYN_ARCHBEH of nd2_24516 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24515 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24515;

architecture SYN_ARCHBEH of nd2_24515 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24514 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24514;

architecture SYN_ARCHBEH of nd2_24514 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24513 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24513;

architecture SYN_ARCHBEH of nd2_24513 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24512 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24512;

architecture SYN_ARCHBEH of nd2_24512 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24511 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24511;

architecture SYN_ARCHBEH of nd2_24511 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24510 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24510;

architecture SYN_ARCHBEH of nd2_24510 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24509 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24509;

architecture SYN_ARCHBEH of nd2_24509 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24508 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24508;

architecture SYN_ARCHBEH of nd2_24508 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24507 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24507;

architecture SYN_ARCHBEH of nd2_24507 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24506 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24506;

architecture SYN_ARCHBEH of nd2_24506 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24505 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24505;

architecture SYN_ARCHBEH of nd2_24505 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24504 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24504;

architecture SYN_ARCHBEH of nd2_24504 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24503 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24503;

architecture SYN_ARCHBEH of nd2_24503 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24502 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24502;

architecture SYN_ARCHBEH of nd2_24502 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24501 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24501;

architecture SYN_ARCHBEH of nd2_24501 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24500 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24500;

architecture SYN_ARCHBEH of nd2_24500 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24499 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24499;

architecture SYN_ARCHBEH of nd2_24499 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24498 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24498;

architecture SYN_ARCHBEH of nd2_24498 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24497 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24497;

architecture SYN_ARCHBEH of nd2_24497 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24496 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24496;

architecture SYN_ARCHBEH of nd2_24496 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24495 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24495;

architecture SYN_ARCHBEH of nd2_24495 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24494 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24494;

architecture SYN_ARCHBEH of nd2_24494 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24493 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24493;

architecture SYN_ARCHBEH of nd2_24493 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24492 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24492;

architecture SYN_ARCHBEH of nd2_24492 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24491 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24491;

architecture SYN_ARCHBEH of nd2_24491 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24490 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24490;

architecture SYN_ARCHBEH of nd2_24490 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24489 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24489;

architecture SYN_ARCHBEH of nd2_24489 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24488 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24488;

architecture SYN_ARCHBEH of nd2_24488 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24487 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24487;

architecture SYN_ARCHBEH of nd2_24487 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24486 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24486;

architecture SYN_ARCHBEH of nd2_24486 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24485 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24485;

architecture SYN_ARCHBEH of nd2_24485 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24484 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24484;

architecture SYN_ARCHBEH of nd2_24484 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24483 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24483;

architecture SYN_ARCHBEH of nd2_24483 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24482 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24482;

architecture SYN_ARCHBEH of nd2_24482 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24481 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24481;

architecture SYN_ARCHBEH of nd2_24481 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24480 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24480;

architecture SYN_ARCHBEH of nd2_24480 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24479 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24479;

architecture SYN_ARCHBEH of nd2_24479 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24478 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24478;

architecture SYN_ARCHBEH of nd2_24478 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24477 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24477;

architecture SYN_ARCHBEH of nd2_24477 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24476 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24476;

architecture SYN_ARCHBEH of nd2_24476 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24475 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24475;

architecture SYN_ARCHBEH of nd2_24475 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24474 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24474;

architecture SYN_ARCHBEH of nd2_24474 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24473 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24473;

architecture SYN_ARCHBEH of nd2_24473 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24472 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24472;

architecture SYN_ARCHBEH of nd2_24472 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24471 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24471;

architecture SYN_ARCHBEH of nd2_24471 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24470 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24470;

architecture SYN_ARCHBEH of nd2_24470 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24469 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24469;

architecture SYN_ARCHBEH of nd2_24469 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24468 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24468;

architecture SYN_ARCHBEH of nd2_24468 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24467 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24467;

architecture SYN_ARCHBEH of nd2_24467 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24466 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24466;

architecture SYN_ARCHBEH of nd2_24466 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24465 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24465;

architecture SYN_ARCHBEH of nd2_24465 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24464 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24464;

architecture SYN_ARCHBEH of nd2_24464 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24463 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24463;

architecture SYN_ARCHBEH of nd2_24463 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24462 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24462;

architecture SYN_ARCHBEH of nd2_24462 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24461 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24461;

architecture SYN_ARCHBEH of nd2_24461 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24460 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24460;

architecture SYN_ARCHBEH of nd2_24460 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24459 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24459;

architecture SYN_ARCHBEH of nd2_24459 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24458 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24458;

architecture SYN_ARCHBEH of nd2_24458 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24457 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24457;

architecture SYN_ARCHBEH of nd2_24457 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24456 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24456;

architecture SYN_ARCHBEH of nd2_24456 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24455 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24455;

architecture SYN_ARCHBEH of nd2_24455 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24454 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24454;

architecture SYN_ARCHBEH of nd2_24454 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24453 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24453;

architecture SYN_ARCHBEH of nd2_24453 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24452 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24452;

architecture SYN_ARCHBEH of nd2_24452 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24451 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24451;

architecture SYN_ARCHBEH of nd2_24451 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24450 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24450;

architecture SYN_ARCHBEH of nd2_24450 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24449 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24449;

architecture SYN_ARCHBEH of nd2_24449 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24448 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24448;

architecture SYN_ARCHBEH of nd2_24448 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24447 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24447;

architecture SYN_ARCHBEH of nd2_24447 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24446 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24446;

architecture SYN_ARCHBEH of nd2_24446 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24445 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24445;

architecture SYN_ARCHBEH of nd2_24445 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24444 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24444;

architecture SYN_ARCHBEH of nd2_24444 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24443 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24443;

architecture SYN_ARCHBEH of nd2_24443 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24442 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24442;

architecture SYN_ARCHBEH of nd2_24442 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24441 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24441;

architecture SYN_ARCHBEH of nd2_24441 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24440 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24440;

architecture SYN_ARCHBEH of nd2_24440 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24439 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24439;

architecture SYN_ARCHBEH of nd2_24439 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24438 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24438;

architecture SYN_ARCHBEH of nd2_24438 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24437 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24437;

architecture SYN_ARCHBEH of nd2_24437 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24436 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24436;

architecture SYN_ARCHBEH of nd2_24436 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24435 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24435;

architecture SYN_ARCHBEH of nd2_24435 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24434 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24434;

architecture SYN_ARCHBEH of nd2_24434 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24433 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24433;

architecture SYN_ARCHBEH of nd2_24433 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24432 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24432;

architecture SYN_ARCHBEH of nd2_24432 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24431 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24431;

architecture SYN_ARCHBEH of nd2_24431 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24430 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24430;

architecture SYN_ARCHBEH of nd2_24430 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24429 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24429;

architecture SYN_ARCHBEH of nd2_24429 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24428 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24428;

architecture SYN_ARCHBEH of nd2_24428 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24427 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24427;

architecture SYN_ARCHBEH of nd2_24427 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24426 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24426;

architecture SYN_ARCHBEH of nd2_24426 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24425 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24425;

architecture SYN_ARCHBEH of nd2_24425 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24424 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24424;

architecture SYN_ARCHBEH of nd2_24424 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24423 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24423;

architecture SYN_ARCHBEH of nd2_24423 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24422 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24422;

architecture SYN_ARCHBEH of nd2_24422 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24421 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24421;

architecture SYN_ARCHBEH of nd2_24421 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24420 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24420;

architecture SYN_ARCHBEH of nd2_24420 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24419 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24419;

architecture SYN_ARCHBEH of nd2_24419 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24418 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24418;

architecture SYN_ARCHBEH of nd2_24418 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24417 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24417;

architecture SYN_ARCHBEH of nd2_24417 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24416 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24416;

architecture SYN_ARCHBEH of nd2_24416 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24415 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24415;

architecture SYN_ARCHBEH of nd2_24415 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24414 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24414;

architecture SYN_ARCHBEH of nd2_24414 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24413 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24413;

architecture SYN_ARCHBEH of nd2_24413 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24412 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24412;

architecture SYN_ARCHBEH of nd2_24412 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24411 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24411;

architecture SYN_ARCHBEH of nd2_24411 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24410 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24410;

architecture SYN_ARCHBEH of nd2_24410 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24409 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24409;

architecture SYN_ARCHBEH of nd2_24409 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24408 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24408;

architecture SYN_ARCHBEH of nd2_24408 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24407 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24407;

architecture SYN_ARCHBEH of nd2_24407 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24406 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24406;

architecture SYN_ARCHBEH of nd2_24406 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24405 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24405;

architecture SYN_ARCHBEH of nd2_24405 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24404 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24404;

architecture SYN_ARCHBEH of nd2_24404 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24403 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24403;

architecture SYN_ARCHBEH of nd2_24403 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24402 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24402;

architecture SYN_ARCHBEH of nd2_24402 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24401 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24401;

architecture SYN_ARCHBEH of nd2_24401 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24400 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24400;

architecture SYN_ARCHBEH of nd2_24400 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24399 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24399;

architecture SYN_ARCHBEH of nd2_24399 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24398 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24398;

architecture SYN_ARCHBEH of nd2_24398 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24397 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24397;

architecture SYN_ARCHBEH of nd2_24397 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24396 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24396;

architecture SYN_ARCHBEH of nd2_24396 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24395 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24395;

architecture SYN_ARCHBEH of nd2_24395 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24394 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24394;

architecture SYN_ARCHBEH of nd2_24394 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24393 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24393;

architecture SYN_ARCHBEH of nd2_24393 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24392 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24392;

architecture SYN_ARCHBEH of nd2_24392 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24391 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24391;

architecture SYN_ARCHBEH of nd2_24391 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24390 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24390;

architecture SYN_ARCHBEH of nd2_24390 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24389 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24389;

architecture SYN_ARCHBEH of nd2_24389 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24388 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24388;

architecture SYN_ARCHBEH of nd2_24388 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24387 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24387;

architecture SYN_ARCHBEH of nd2_24387 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24386 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24386;

architecture SYN_ARCHBEH of nd2_24386 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24385 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24385;

architecture SYN_ARCHBEH of nd2_24385 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8623 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8623;

architecture SYN_ARCHSTRUCT of iv_8623 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8622 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8622;

architecture SYN_ARCHSTRUCT of iv_8622 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8621 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8621;

architecture SYN_ARCHSTRUCT of iv_8621 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8620 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8620;

architecture SYN_ARCHSTRUCT of iv_8620 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8619 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8619;

architecture SYN_ARCHSTRUCT of iv_8619 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8618 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8618;

architecture SYN_ARCHSTRUCT of iv_8618 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8617 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8617;

architecture SYN_ARCHSTRUCT of iv_8617 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8616 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8616;

architecture SYN_ARCHSTRUCT of iv_8616 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8615 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8615;

architecture SYN_ARCHSTRUCT of iv_8615 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8614 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8614;

architecture SYN_ARCHSTRUCT of iv_8614 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8613 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8613;

architecture SYN_ARCHSTRUCT of iv_8613 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8612 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8612;

architecture SYN_ARCHSTRUCT of iv_8612 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8611 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8611;

architecture SYN_ARCHSTRUCT of iv_8611 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8610 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8610;

architecture SYN_ARCHSTRUCT of iv_8610 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8609 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8609;

architecture SYN_ARCHSTRUCT of iv_8609 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8608 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8608;

architecture SYN_ARCHSTRUCT of iv_8608 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8607 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8607;

architecture SYN_ARCHSTRUCT of iv_8607 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8606 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8606;

architecture SYN_ARCHSTRUCT of iv_8606 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8605 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8605;

architecture SYN_ARCHSTRUCT of iv_8605 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8604 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8604;

architecture SYN_ARCHSTRUCT of iv_8604 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8603 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8603;

architecture SYN_ARCHSTRUCT of iv_8603 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8602 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8602;

architecture SYN_ARCHSTRUCT of iv_8602 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8601 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8601;

architecture SYN_ARCHSTRUCT of iv_8601 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8600 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8600;

architecture SYN_ARCHSTRUCT of iv_8600 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8599 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8599;

architecture SYN_ARCHSTRUCT of iv_8599 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8598 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8598;

architecture SYN_ARCHSTRUCT of iv_8598 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8597 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8597;

architecture SYN_ARCHSTRUCT of iv_8597 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8596 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8596;

architecture SYN_ARCHSTRUCT of iv_8596 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8595 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8595;

architecture SYN_ARCHSTRUCT of iv_8595 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8594 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8594;

architecture SYN_ARCHSTRUCT of iv_8594 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8593 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8593;

architecture SYN_ARCHSTRUCT of iv_8593 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8592 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8592;

architecture SYN_ARCHSTRUCT of iv_8592 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8591 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8591;

architecture SYN_ARCHSTRUCT of iv_8591 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8590 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8590;

architecture SYN_ARCHSTRUCT of iv_8590 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8589 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8589;

architecture SYN_ARCHSTRUCT of iv_8589 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8588 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8588;

architecture SYN_ARCHSTRUCT of iv_8588 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8587 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8587;

architecture SYN_ARCHSTRUCT of iv_8587 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8586 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8586;

architecture SYN_ARCHSTRUCT of iv_8586 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8585 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8585;

architecture SYN_ARCHSTRUCT of iv_8585 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8584 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8584;

architecture SYN_ARCHSTRUCT of iv_8584 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8583 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8583;

architecture SYN_ARCHSTRUCT of iv_8583 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8582 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8582;

architecture SYN_ARCHSTRUCT of iv_8582 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8581 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8581;

architecture SYN_ARCHSTRUCT of iv_8581 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8580 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8580;

architecture SYN_ARCHSTRUCT of iv_8580 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8579 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8579;

architecture SYN_ARCHSTRUCT of iv_8579 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8578 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8578;

architecture SYN_ARCHSTRUCT of iv_8578 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8577 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8577;

architecture SYN_ARCHSTRUCT of iv_8577 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8576 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8576;

architecture SYN_ARCHSTRUCT of iv_8576 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8575 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8575;

architecture SYN_ARCHSTRUCT of iv_8575 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8574 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8574;

architecture SYN_ARCHSTRUCT of iv_8574 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8573 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8573;

architecture SYN_ARCHSTRUCT of iv_8573 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8572 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8572;

architecture SYN_ARCHSTRUCT of iv_8572 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8571 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8571;

architecture SYN_ARCHSTRUCT of iv_8571 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8570 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8570;

architecture SYN_ARCHSTRUCT of iv_8570 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8569 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8569;

architecture SYN_ARCHSTRUCT of iv_8569 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8568 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8568;

architecture SYN_ARCHSTRUCT of iv_8568 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8567 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8567;

architecture SYN_ARCHSTRUCT of iv_8567 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8566 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8566;

architecture SYN_ARCHSTRUCT of iv_8566 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8565 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8565;

architecture SYN_ARCHSTRUCT of iv_8565 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8564 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8564;

architecture SYN_ARCHSTRUCT of iv_8564 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8563 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8563;

architecture SYN_ARCHSTRUCT of iv_8563 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8562 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8562;

architecture SYN_ARCHSTRUCT of iv_8562 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8561 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8561;

architecture SYN_ARCHSTRUCT of iv_8561 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8560 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8560;

architecture SYN_ARCHSTRUCT of iv_8560 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8559 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8559;

architecture SYN_ARCHSTRUCT of iv_8559 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8558 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8558;

architecture SYN_ARCHSTRUCT of iv_8558 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8557 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8557;

architecture SYN_ARCHSTRUCT of iv_8557 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8556 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8556;

architecture SYN_ARCHSTRUCT of iv_8556 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8555 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8555;

architecture SYN_ARCHSTRUCT of iv_8555 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8554 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8554;

architecture SYN_ARCHSTRUCT of iv_8554 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8553 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8553;

architecture SYN_ARCHSTRUCT of iv_8553 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8552 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8552;

architecture SYN_ARCHSTRUCT of iv_8552 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8551 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8551;

architecture SYN_ARCHSTRUCT of iv_8551 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8550 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8550;

architecture SYN_ARCHSTRUCT of iv_8550 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8549 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8549;

architecture SYN_ARCHSTRUCT of iv_8549 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8548 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8548;

architecture SYN_ARCHSTRUCT of iv_8548 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8547 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8547;

architecture SYN_ARCHSTRUCT of iv_8547 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8546 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8546;

architecture SYN_ARCHSTRUCT of iv_8546 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8545 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8545;

architecture SYN_ARCHSTRUCT of iv_8545 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8544 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8544;

architecture SYN_ARCHSTRUCT of iv_8544 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8543 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8543;

architecture SYN_ARCHSTRUCT of iv_8543 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8542 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8542;

architecture SYN_ARCHSTRUCT of iv_8542 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8541 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8541;

architecture SYN_ARCHSTRUCT of iv_8541 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8540 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8540;

architecture SYN_ARCHSTRUCT of iv_8540 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8539 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8539;

architecture SYN_ARCHSTRUCT of iv_8539 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8538 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8538;

architecture SYN_ARCHSTRUCT of iv_8538 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8537 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8537;

architecture SYN_ARCHSTRUCT of iv_8537 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8536 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8536;

architecture SYN_ARCHSTRUCT of iv_8536 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8535 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8535;

architecture SYN_ARCHSTRUCT of iv_8535 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8534 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8534;

architecture SYN_ARCHSTRUCT of iv_8534 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8533 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8533;

architecture SYN_ARCHSTRUCT of iv_8533 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8532 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8532;

architecture SYN_ARCHSTRUCT of iv_8532 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8531 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8531;

architecture SYN_ARCHSTRUCT of iv_8531 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8530 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8530;

architecture SYN_ARCHSTRUCT of iv_8530 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8529 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8529;

architecture SYN_ARCHSTRUCT of iv_8529 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8528 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8528;

architecture SYN_ARCHSTRUCT of iv_8528 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8527 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8527;

architecture SYN_ARCHSTRUCT of iv_8527 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8526 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8526;

architecture SYN_ARCHSTRUCT of iv_8526 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8525 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8525;

architecture SYN_ARCHSTRUCT of iv_8525 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8524 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8524;

architecture SYN_ARCHSTRUCT of iv_8524 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8523 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8523;

architecture SYN_ARCHSTRUCT of iv_8523 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8522 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8522;

architecture SYN_ARCHSTRUCT of iv_8522 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8521 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8521;

architecture SYN_ARCHSTRUCT of iv_8521 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8520 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8520;

architecture SYN_ARCHSTRUCT of iv_8520 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8519 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8519;

architecture SYN_ARCHSTRUCT of iv_8519 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8518 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8518;

architecture SYN_ARCHSTRUCT of iv_8518 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8517 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8517;

architecture SYN_ARCHSTRUCT of iv_8517 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8516 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8516;

architecture SYN_ARCHSTRUCT of iv_8516 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8515 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8515;

architecture SYN_ARCHSTRUCT of iv_8515 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8514 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8514;

architecture SYN_ARCHSTRUCT of iv_8514 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8513 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8513;

architecture SYN_ARCHSTRUCT of iv_8513 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8512 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8512;

architecture SYN_ARCHSTRUCT of iv_8512 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8511 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8511;

architecture SYN_ARCHSTRUCT of iv_8511 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8510 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8510;

architecture SYN_ARCHSTRUCT of iv_8510 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8509 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8509;

architecture SYN_ARCHSTRUCT of iv_8509 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8508 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8508;

architecture SYN_ARCHSTRUCT of iv_8508 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8507 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8507;

architecture SYN_ARCHSTRUCT of iv_8507 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8506 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8506;

architecture SYN_ARCHSTRUCT of iv_8506 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8505 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8505;

architecture SYN_ARCHSTRUCT of iv_8505 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8504 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8504;

architecture SYN_ARCHSTRUCT of iv_8504 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8503 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8503;

architecture SYN_ARCHSTRUCT of iv_8503 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8502 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8502;

architecture SYN_ARCHSTRUCT of iv_8502 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8501 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8501;

architecture SYN_ARCHSTRUCT of iv_8501 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8500 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8500;

architecture SYN_ARCHSTRUCT of iv_8500 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8499 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8499;

architecture SYN_ARCHSTRUCT of iv_8499 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8498 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8498;

architecture SYN_ARCHSTRUCT of iv_8498 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8497 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8497;

architecture SYN_ARCHSTRUCT of iv_8497 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8496 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8496;

architecture SYN_ARCHSTRUCT of iv_8496 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8495 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8495;

architecture SYN_ARCHSTRUCT of iv_8495 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8494 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8494;

architecture SYN_ARCHSTRUCT of iv_8494 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8493 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8493;

architecture SYN_ARCHSTRUCT of iv_8493 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8492 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8492;

architecture SYN_ARCHSTRUCT of iv_8492 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8491 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8491;

architecture SYN_ARCHSTRUCT of iv_8491 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8490 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8490;

architecture SYN_ARCHSTRUCT of iv_8490 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8489 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8489;

architecture SYN_ARCHSTRUCT of iv_8489 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8488 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8488;

architecture SYN_ARCHSTRUCT of iv_8488 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8487 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8487;

architecture SYN_ARCHSTRUCT of iv_8487 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8486 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8486;

architecture SYN_ARCHSTRUCT of iv_8486 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8485 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8485;

architecture SYN_ARCHSTRUCT of iv_8485 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8484 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8484;

architecture SYN_ARCHSTRUCT of iv_8484 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8483 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8483;

architecture SYN_ARCHSTRUCT of iv_8483 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8482 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8482;

architecture SYN_ARCHSTRUCT of iv_8482 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8481 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8481;

architecture SYN_ARCHSTRUCT of iv_8481 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8480 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8480;

architecture SYN_ARCHSTRUCT of iv_8480 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8479 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8479;

architecture SYN_ARCHSTRUCT of iv_8479 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8478 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8478;

architecture SYN_ARCHSTRUCT of iv_8478 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8477 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8477;

architecture SYN_ARCHSTRUCT of iv_8477 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8476 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8476;

architecture SYN_ARCHSTRUCT of iv_8476 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8475 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8475;

architecture SYN_ARCHSTRUCT of iv_8475 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8474 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8474;

architecture SYN_ARCHSTRUCT of iv_8474 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8473 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8473;

architecture SYN_ARCHSTRUCT of iv_8473 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8472 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8472;

architecture SYN_ARCHSTRUCT of iv_8472 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8471 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8471;

architecture SYN_ARCHSTRUCT of iv_8471 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8470 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8470;

architecture SYN_ARCHSTRUCT of iv_8470 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8469 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8469;

architecture SYN_ARCHSTRUCT of iv_8469 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8468 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8468;

architecture SYN_ARCHSTRUCT of iv_8468 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8467 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8467;

architecture SYN_ARCHSTRUCT of iv_8467 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8466 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8466;

architecture SYN_ARCHSTRUCT of iv_8466 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8465 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8465;

architecture SYN_ARCHSTRUCT of iv_8465 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8464 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8464;

architecture SYN_ARCHSTRUCT of iv_8464 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8463 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8463;

architecture SYN_ARCHSTRUCT of iv_8463 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8462 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8462;

architecture SYN_ARCHSTRUCT of iv_8462 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8461 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8461;

architecture SYN_ARCHSTRUCT of iv_8461 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8460 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8460;

architecture SYN_ARCHSTRUCT of iv_8460 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8459 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8459;

architecture SYN_ARCHSTRUCT of iv_8459 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8458 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8458;

architecture SYN_ARCHSTRUCT of iv_8458 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8457 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8457;

architecture SYN_ARCHSTRUCT of iv_8457 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8456 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8456;

architecture SYN_ARCHSTRUCT of iv_8456 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8455 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8455;

architecture SYN_ARCHSTRUCT of iv_8455 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8454 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8454;

architecture SYN_ARCHSTRUCT of iv_8454 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8453 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8453;

architecture SYN_ARCHSTRUCT of iv_8453 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8452 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8452;

architecture SYN_ARCHSTRUCT of iv_8452 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8451 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8451;

architecture SYN_ARCHSTRUCT of iv_8451 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8450 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8450;

architecture SYN_ARCHSTRUCT of iv_8450 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8449 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8449;

architecture SYN_ARCHSTRUCT of iv_8449 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8448 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8448;

architecture SYN_ARCHSTRUCT of iv_8448 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8447 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8447;

architecture SYN_ARCHSTRUCT of iv_8447 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8446 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8446;

architecture SYN_ARCHSTRUCT of iv_8446 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8445 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8445;

architecture SYN_ARCHSTRUCT of iv_8445 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8444 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8444;

architecture SYN_ARCHSTRUCT of iv_8444 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8443 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8443;

architecture SYN_ARCHSTRUCT of iv_8443 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8442 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8442;

architecture SYN_ARCHSTRUCT of iv_8442 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8441 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8441;

architecture SYN_ARCHSTRUCT of iv_8441 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8440 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8440;

architecture SYN_ARCHSTRUCT of iv_8440 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8439 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8439;

architecture SYN_ARCHSTRUCT of iv_8439 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8438 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8438;

architecture SYN_ARCHSTRUCT of iv_8438 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8437 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8437;

architecture SYN_ARCHSTRUCT of iv_8437 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8436 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8436;

architecture SYN_ARCHSTRUCT of iv_8436 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8435 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8435;

architecture SYN_ARCHSTRUCT of iv_8435 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8434 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8434;

architecture SYN_ARCHSTRUCT of iv_8434 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8433 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8433;

architecture SYN_ARCHSTRUCT of iv_8433 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8432 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8432;

architecture SYN_ARCHSTRUCT of iv_8432 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8431 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8431;

architecture SYN_ARCHSTRUCT of iv_8431 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8430 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8430;

architecture SYN_ARCHSTRUCT of iv_8430 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8429 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8429;

architecture SYN_ARCHSTRUCT of iv_8429 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8428 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8428;

architecture SYN_ARCHSTRUCT of iv_8428 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8427 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8427;

architecture SYN_ARCHSTRUCT of iv_8427 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8426 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8426;

architecture SYN_ARCHSTRUCT of iv_8426 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8425 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8425;

architecture SYN_ARCHSTRUCT of iv_8425 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8424 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8424;

architecture SYN_ARCHSTRUCT of iv_8424 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8423 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8423;

architecture SYN_ARCHSTRUCT of iv_8423 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8422 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8422;

architecture SYN_ARCHSTRUCT of iv_8422 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8421 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8421;

architecture SYN_ARCHSTRUCT of iv_8421 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8420 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8420;

architecture SYN_ARCHSTRUCT of iv_8420 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8419 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8419;

architecture SYN_ARCHSTRUCT of iv_8419 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8418 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8418;

architecture SYN_ARCHSTRUCT of iv_8418 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8417 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8417;

architecture SYN_ARCHSTRUCT of iv_8417 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8416 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8416;

architecture SYN_ARCHSTRUCT of iv_8416 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8415 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8415;

architecture SYN_ARCHSTRUCT of iv_8415 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8414 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8414;

architecture SYN_ARCHSTRUCT of iv_8414 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8413 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8413;

architecture SYN_ARCHSTRUCT of iv_8413 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8412 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8412;

architecture SYN_ARCHSTRUCT of iv_8412 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8411 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8411;

architecture SYN_ARCHSTRUCT of iv_8411 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8410 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8410;

architecture SYN_ARCHSTRUCT of iv_8410 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8409 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8409;

architecture SYN_ARCHSTRUCT of iv_8409 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8408 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8408;

architecture SYN_ARCHSTRUCT of iv_8408 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8407 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8407;

architecture SYN_ARCHSTRUCT of iv_8407 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8406 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8406;

architecture SYN_ARCHSTRUCT of iv_8406 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8405 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8405;

architecture SYN_ARCHSTRUCT of iv_8405 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8404 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8404;

architecture SYN_ARCHSTRUCT of iv_8404 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8403 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8403;

architecture SYN_ARCHSTRUCT of iv_8403 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8402 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8402;

architecture SYN_ARCHSTRUCT of iv_8402 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8401 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8401;

architecture SYN_ARCHSTRUCT of iv_8401 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8400 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8400;

architecture SYN_ARCHSTRUCT of iv_8400 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8399 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8399;

architecture SYN_ARCHSTRUCT of iv_8399 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8398 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8398;

architecture SYN_ARCHSTRUCT of iv_8398 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8397 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8397;

architecture SYN_ARCHSTRUCT of iv_8397 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8396 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8396;

architecture SYN_ARCHSTRUCT of iv_8396 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8395 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8395;

architecture SYN_ARCHSTRUCT of iv_8395 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8394 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8394;

architecture SYN_ARCHSTRUCT of iv_8394 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8393 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8393;

architecture SYN_ARCHSTRUCT of iv_8393 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8392 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8392;

architecture SYN_ARCHSTRUCT of iv_8392 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8391 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8391;

architecture SYN_ARCHSTRUCT of iv_8391 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8390 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8390;

architecture SYN_ARCHSTRUCT of iv_8390 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8389 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8389;

architecture SYN_ARCHSTRUCT of iv_8389 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8388 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8388;

architecture SYN_ARCHSTRUCT of iv_8388 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8387 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8387;

architecture SYN_ARCHSTRUCT of iv_8387 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8386 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8386;

architecture SYN_ARCHSTRUCT of iv_8386 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8385 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8385;

architecture SYN_ARCHSTRUCT of iv_8385 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8384 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8384;

architecture SYN_ARCHSTRUCT of iv_8384 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8383 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8383;

architecture SYN_ARCHSTRUCT of iv_8383 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8382 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8382;

architecture SYN_ARCHSTRUCT of iv_8382 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8381 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8381;

architecture SYN_ARCHSTRUCT of iv_8381 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8380 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8380;

architecture SYN_ARCHSTRUCT of iv_8380 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8379 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8379;

architecture SYN_ARCHSTRUCT of iv_8379 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8378 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8378;

architecture SYN_ARCHSTRUCT of iv_8378 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8377 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8377;

architecture SYN_ARCHSTRUCT of iv_8377 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8376 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8376;

architecture SYN_ARCHSTRUCT of iv_8376 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8375 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8375;

architecture SYN_ARCHSTRUCT of iv_8375 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8374 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8374;

architecture SYN_ARCHSTRUCT of iv_8374 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8373 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8373;

architecture SYN_ARCHSTRUCT of iv_8373 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8372 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8372;

architecture SYN_ARCHSTRUCT of iv_8372 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8371 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8371;

architecture SYN_ARCHSTRUCT of iv_8371 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8370 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8370;

architecture SYN_ARCHSTRUCT of iv_8370 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8369 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8369;

architecture SYN_ARCHSTRUCT of iv_8369 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8368 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8368;

architecture SYN_ARCHSTRUCT of iv_8368 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8367 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8367;

architecture SYN_ARCHSTRUCT of iv_8367 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8366 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8366;

architecture SYN_ARCHSTRUCT of iv_8366 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8365 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8365;

architecture SYN_ARCHSTRUCT of iv_8365 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8364 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8364;

architecture SYN_ARCHSTRUCT of iv_8364 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8363 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8363;

architecture SYN_ARCHSTRUCT of iv_8363 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8362 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8362;

architecture SYN_ARCHSTRUCT of iv_8362 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8361 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8361;

architecture SYN_ARCHSTRUCT of iv_8361 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8360 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8360;

architecture SYN_ARCHSTRUCT of iv_8360 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8359 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8359;

architecture SYN_ARCHSTRUCT of iv_8359 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8358 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8358;

architecture SYN_ARCHSTRUCT of iv_8358 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8357 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8357;

architecture SYN_ARCHSTRUCT of iv_8357 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8356 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8356;

architecture SYN_ARCHSTRUCT of iv_8356 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8355 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8355;

architecture SYN_ARCHSTRUCT of iv_8355 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8354 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8354;

architecture SYN_ARCHSTRUCT of iv_8354 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8353 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8353;

architecture SYN_ARCHSTRUCT of iv_8353 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8352 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8352;

architecture SYN_ARCHSTRUCT of iv_8352 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8351 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8351;

architecture SYN_ARCHSTRUCT of iv_8351 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8350 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8350;

architecture SYN_ARCHSTRUCT of iv_8350 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8349 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8349;

architecture SYN_ARCHSTRUCT of iv_8349 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8348 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8348;

architecture SYN_ARCHSTRUCT of iv_8348 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8347 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8347;

architecture SYN_ARCHSTRUCT of iv_8347 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8346 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8346;

architecture SYN_ARCHSTRUCT of iv_8346 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8345 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8345;

architecture SYN_ARCHSTRUCT of iv_8345 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8344 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8344;

architecture SYN_ARCHSTRUCT of iv_8344 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8343 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8343;

architecture SYN_ARCHSTRUCT of iv_8343 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8342 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8342;

architecture SYN_ARCHSTRUCT of iv_8342 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8341 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8341;

architecture SYN_ARCHSTRUCT of iv_8341 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8340 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8340;

architecture SYN_ARCHSTRUCT of iv_8340 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8339 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8339;

architecture SYN_ARCHSTRUCT of iv_8339 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8338 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8338;

architecture SYN_ARCHSTRUCT of iv_8338 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8337 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8337;

architecture SYN_ARCHSTRUCT of iv_8337 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8336 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8336;

architecture SYN_ARCHSTRUCT of iv_8336 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8335 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8335;

architecture SYN_ARCHSTRUCT of iv_8335 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8334 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8334;

architecture SYN_ARCHSTRUCT of iv_8334 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8333 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8333;

architecture SYN_ARCHSTRUCT of iv_8333 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8332 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8332;

architecture SYN_ARCHSTRUCT of iv_8332 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8331 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8331;

architecture SYN_ARCHSTRUCT of iv_8331 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8330 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8330;

architecture SYN_ARCHSTRUCT of iv_8330 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8329 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8329;

architecture SYN_ARCHSTRUCT of iv_8329 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8328 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8328;

architecture SYN_ARCHSTRUCT of iv_8328 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8327 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8327;

architecture SYN_ARCHSTRUCT of iv_8327 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8326 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8326;

architecture SYN_ARCHSTRUCT of iv_8326 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8325 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8325;

architecture SYN_ARCHSTRUCT of iv_8325 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8324 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8324;

architecture SYN_ARCHSTRUCT of iv_8324 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8323 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8323;

architecture SYN_ARCHSTRUCT of iv_8323 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8322 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8322;

architecture SYN_ARCHSTRUCT of iv_8322 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8321 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8321;

architecture SYN_ARCHSTRUCT of iv_8321 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8320 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8320;

architecture SYN_ARCHSTRUCT of iv_8320 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8319 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8319;

architecture SYN_ARCHSTRUCT of iv_8319 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8318 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8318;

architecture SYN_ARCHSTRUCT of iv_8318 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8317 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8317;

architecture SYN_ARCHSTRUCT of iv_8317 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8316 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8316;

architecture SYN_ARCHSTRUCT of iv_8316 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8315 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8315;

architecture SYN_ARCHSTRUCT of iv_8315 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8314 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8314;

architecture SYN_ARCHSTRUCT of iv_8314 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8313 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8313;

architecture SYN_ARCHSTRUCT of iv_8313 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8312 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8312;

architecture SYN_ARCHSTRUCT of iv_8312 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8311 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8311;

architecture SYN_ARCHSTRUCT of iv_8311 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8310 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8310;

architecture SYN_ARCHSTRUCT of iv_8310 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8309 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8309;

architecture SYN_ARCHSTRUCT of iv_8309 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8308 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8308;

architecture SYN_ARCHSTRUCT of iv_8308 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8307 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8307;

architecture SYN_ARCHSTRUCT of iv_8307 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8306 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8306;

architecture SYN_ARCHSTRUCT of iv_8306 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8305 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8305;

architecture SYN_ARCHSTRUCT of iv_8305 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8304 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8304;

architecture SYN_ARCHSTRUCT of iv_8304 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8303 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8303;

architecture SYN_ARCHSTRUCT of iv_8303 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8302 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8302;

architecture SYN_ARCHSTRUCT of iv_8302 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8301 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8301;

architecture SYN_ARCHSTRUCT of iv_8301 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8300 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8300;

architecture SYN_ARCHSTRUCT of iv_8300 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8299 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8299;

architecture SYN_ARCHSTRUCT of iv_8299 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8298 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8298;

architecture SYN_ARCHSTRUCT of iv_8298 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8297 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8297;

architecture SYN_ARCHSTRUCT of iv_8297 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8296 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8296;

architecture SYN_ARCHSTRUCT of iv_8296 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8295 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8295;

architecture SYN_ARCHSTRUCT of iv_8295 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8294 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8294;

architecture SYN_ARCHSTRUCT of iv_8294 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8293 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8293;

architecture SYN_ARCHSTRUCT of iv_8293 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8292 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8292;

architecture SYN_ARCHSTRUCT of iv_8292 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8291 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8291;

architecture SYN_ARCHSTRUCT of iv_8291 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8290 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8290;

architecture SYN_ARCHSTRUCT of iv_8290 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8289 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8289;

architecture SYN_ARCHSTRUCT of iv_8289 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8288 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8288;

architecture SYN_ARCHSTRUCT of iv_8288 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8287 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8287;

architecture SYN_ARCHSTRUCT of iv_8287 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8286 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8286;

architecture SYN_ARCHSTRUCT of iv_8286 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8285 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8285;

architecture SYN_ARCHSTRUCT of iv_8285 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8284 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8284;

architecture SYN_ARCHSTRUCT of iv_8284 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8283 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8283;

architecture SYN_ARCHSTRUCT of iv_8283 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8282 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8282;

architecture SYN_ARCHSTRUCT of iv_8282 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8281 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8281;

architecture SYN_ARCHSTRUCT of iv_8281 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8280 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8280;

architecture SYN_ARCHSTRUCT of iv_8280 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8279 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8279;

architecture SYN_ARCHSTRUCT of iv_8279 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8278 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8278;

architecture SYN_ARCHSTRUCT of iv_8278 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8277 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8277;

architecture SYN_ARCHSTRUCT of iv_8277 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8276 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8276;

architecture SYN_ARCHSTRUCT of iv_8276 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8275 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8275;

architecture SYN_ARCHSTRUCT of iv_8275 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8274 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8274;

architecture SYN_ARCHSTRUCT of iv_8274 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8273 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8273;

architecture SYN_ARCHSTRUCT of iv_8273 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8272 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8272;

architecture SYN_ARCHSTRUCT of iv_8272 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8271 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8271;

architecture SYN_ARCHSTRUCT of iv_8271 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8270 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8270;

architecture SYN_ARCHSTRUCT of iv_8270 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8269 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8269;

architecture SYN_ARCHSTRUCT of iv_8269 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8268 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8268;

architecture SYN_ARCHSTRUCT of iv_8268 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8267 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8267;

architecture SYN_ARCHSTRUCT of iv_8267 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8266 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8266;

architecture SYN_ARCHSTRUCT of iv_8266 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8265 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8265;

architecture SYN_ARCHSTRUCT of iv_8265 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8264 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8264;

architecture SYN_ARCHSTRUCT of iv_8264 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8263 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8263;

architecture SYN_ARCHSTRUCT of iv_8263 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8262 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8262;

architecture SYN_ARCHSTRUCT of iv_8262 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8261 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8261;

architecture SYN_ARCHSTRUCT of iv_8261 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8260 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8260;

architecture SYN_ARCHSTRUCT of iv_8260 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8259 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8259;

architecture SYN_ARCHSTRUCT of iv_8259 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8258 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8258;

architecture SYN_ARCHSTRUCT of iv_8258 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8257 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8257;

architecture SYN_ARCHSTRUCT of iv_8257 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8256 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8256;

architecture SYN_ARCHSTRUCT of iv_8256 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8255 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8255;

architecture SYN_ARCHSTRUCT of iv_8255 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8254 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8254;

architecture SYN_ARCHSTRUCT of iv_8254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8253 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8253;

architecture SYN_ARCHSTRUCT of iv_8253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8252 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8252;

architecture SYN_ARCHSTRUCT of iv_8252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8251 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8251;

architecture SYN_ARCHSTRUCT of iv_8251 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8250 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8250;

architecture SYN_ARCHSTRUCT of iv_8250 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8249 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8249;

architecture SYN_ARCHSTRUCT of iv_8249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8248 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8248;

architecture SYN_ARCHSTRUCT of iv_8248 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8247 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8247;

architecture SYN_ARCHSTRUCT of iv_8247 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8246 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8246;

architecture SYN_ARCHSTRUCT of iv_8246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8245 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8245;

architecture SYN_ARCHSTRUCT of iv_8245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8244 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8244;

architecture SYN_ARCHSTRUCT of iv_8244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8243 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8243;

architecture SYN_ARCHSTRUCT of iv_8243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8242 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8242;

architecture SYN_ARCHSTRUCT of iv_8242 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8241 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8241;

architecture SYN_ARCHSTRUCT of iv_8241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8240 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8240;

architecture SYN_ARCHSTRUCT of iv_8240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8239 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8239;

architecture SYN_ARCHSTRUCT of iv_8239 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8238 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8238;

architecture SYN_ARCHSTRUCT of iv_8238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8237 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8237;

architecture SYN_ARCHSTRUCT of iv_8237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8236 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8236;

architecture SYN_ARCHSTRUCT of iv_8236 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8235 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8235;

architecture SYN_ARCHSTRUCT of iv_8235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8234 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8234;

architecture SYN_ARCHSTRUCT of iv_8234 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8233 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8233;

architecture SYN_ARCHSTRUCT of iv_8233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8232 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8232;

architecture SYN_ARCHSTRUCT of iv_8232 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8231 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8231;

architecture SYN_ARCHSTRUCT of iv_8231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8230 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8230;

architecture SYN_ARCHSTRUCT of iv_8230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8229 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8229;

architecture SYN_ARCHSTRUCT of iv_8229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8228 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8228;

architecture SYN_ARCHSTRUCT of iv_8228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8227 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8227;

architecture SYN_ARCHSTRUCT of iv_8227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8226 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8226;

architecture SYN_ARCHSTRUCT of iv_8226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8225 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8225;

architecture SYN_ARCHSTRUCT of iv_8225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8224 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8224;

architecture SYN_ARCHSTRUCT of iv_8224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8223 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8223;

architecture SYN_ARCHSTRUCT of iv_8223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8222 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8222;

architecture SYN_ARCHSTRUCT of iv_8222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8221 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8221;

architecture SYN_ARCHSTRUCT of iv_8221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8220 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8220;

architecture SYN_ARCHSTRUCT of iv_8220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8219 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8219;

architecture SYN_ARCHSTRUCT of iv_8219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8218 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8218;

architecture SYN_ARCHSTRUCT of iv_8218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8217 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8217;

architecture SYN_ARCHSTRUCT of iv_8217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8216 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8216;

architecture SYN_ARCHSTRUCT of iv_8216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8215 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8215;

architecture SYN_ARCHSTRUCT of iv_8215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8214 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8214;

architecture SYN_ARCHSTRUCT of iv_8214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8213 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8213;

architecture SYN_ARCHSTRUCT of iv_8213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8212 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8212;

architecture SYN_ARCHSTRUCT of iv_8212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8211 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8211;

architecture SYN_ARCHSTRUCT of iv_8211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8210 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8210;

architecture SYN_ARCHSTRUCT of iv_8210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8209 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8209;

architecture SYN_ARCHSTRUCT of iv_8209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8208 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8208;

architecture SYN_ARCHSTRUCT of iv_8208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8207 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8207;

architecture SYN_ARCHSTRUCT of iv_8207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8206 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8206;

architecture SYN_ARCHSTRUCT of iv_8206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8205 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8205;

architecture SYN_ARCHSTRUCT of iv_8205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8204 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8204;

architecture SYN_ARCHSTRUCT of iv_8204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8203 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8203;

architecture SYN_ARCHSTRUCT of iv_8203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8202 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8202;

architecture SYN_ARCHSTRUCT of iv_8202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8201 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8201;

architecture SYN_ARCHSTRUCT of iv_8201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8200 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8200;

architecture SYN_ARCHSTRUCT of iv_8200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8199 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8199;

architecture SYN_ARCHSTRUCT of iv_8199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8198 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8198;

architecture SYN_ARCHSTRUCT of iv_8198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8197 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8197;

architecture SYN_ARCHSTRUCT of iv_8197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8196 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8196;

architecture SYN_ARCHSTRUCT of iv_8196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8195 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8195;

architecture SYN_ARCHSTRUCT of iv_8195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8194 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8194;

architecture SYN_ARCHSTRUCT of iv_8194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8193 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8193;

architecture SYN_ARCHSTRUCT of iv_8193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8192 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8192;

architecture SYN_ARCHSTRUCT of iv_8192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8191 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8191;

architecture SYN_ARCHSTRUCT of iv_8191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8190 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8190;

architecture SYN_ARCHSTRUCT of iv_8190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8189 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8189;

architecture SYN_ARCHSTRUCT of iv_8189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8188 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8188;

architecture SYN_ARCHSTRUCT of iv_8188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8187 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8187;

architecture SYN_ARCHSTRUCT of iv_8187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8186 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8186;

architecture SYN_ARCHSTRUCT of iv_8186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8185 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8185;

architecture SYN_ARCHSTRUCT of iv_8185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8184 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8184;

architecture SYN_ARCHSTRUCT of iv_8184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8183 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8183;

architecture SYN_ARCHSTRUCT of iv_8183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8182 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8182;

architecture SYN_ARCHSTRUCT of iv_8182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8181 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8181;

architecture SYN_ARCHSTRUCT of iv_8181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8180 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8180;

architecture SYN_ARCHSTRUCT of iv_8180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8179 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8179;

architecture SYN_ARCHSTRUCT of iv_8179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8178 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8178;

architecture SYN_ARCHSTRUCT of iv_8178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8177 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8177;

architecture SYN_ARCHSTRUCT of iv_8177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8176 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8176;

architecture SYN_ARCHSTRUCT of iv_8176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8175 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8175;

architecture SYN_ARCHSTRUCT of iv_8175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8174 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8174;

architecture SYN_ARCHSTRUCT of iv_8174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8173 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8173;

architecture SYN_ARCHSTRUCT of iv_8173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8172 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8172;

architecture SYN_ARCHSTRUCT of iv_8172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8171 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8171;

architecture SYN_ARCHSTRUCT of iv_8171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8170 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8170;

architecture SYN_ARCHSTRUCT of iv_8170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8169 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8169;

architecture SYN_ARCHSTRUCT of iv_8169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8168 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8168;

architecture SYN_ARCHSTRUCT of iv_8168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8167 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8167;

architecture SYN_ARCHSTRUCT of iv_8167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8166 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8166;

architecture SYN_ARCHSTRUCT of iv_8166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8165 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8165;

architecture SYN_ARCHSTRUCT of iv_8165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8164 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8164;

architecture SYN_ARCHSTRUCT of iv_8164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8163 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8163;

architecture SYN_ARCHSTRUCT of iv_8163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8162 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8162;

architecture SYN_ARCHSTRUCT of iv_8162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8161 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8161;

architecture SYN_ARCHSTRUCT of iv_8161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8160 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8160;

architecture SYN_ARCHSTRUCT of iv_8160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8159 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8159;

architecture SYN_ARCHSTRUCT of iv_8159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8158 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8158;

architecture SYN_ARCHSTRUCT of iv_8158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8157 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8157;

architecture SYN_ARCHSTRUCT of iv_8157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8156 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8156;

architecture SYN_ARCHSTRUCT of iv_8156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8155 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8155;

architecture SYN_ARCHSTRUCT of iv_8155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8154 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8154;

architecture SYN_ARCHSTRUCT of iv_8154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8153 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8153;

architecture SYN_ARCHSTRUCT of iv_8153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8152 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8152;

architecture SYN_ARCHSTRUCT of iv_8152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8151 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8151;

architecture SYN_ARCHSTRUCT of iv_8151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8150 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8150;

architecture SYN_ARCHSTRUCT of iv_8150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8149 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8149;

architecture SYN_ARCHSTRUCT of iv_8149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8148 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8148;

architecture SYN_ARCHSTRUCT of iv_8148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8147 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8147;

architecture SYN_ARCHSTRUCT of iv_8147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8146 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8146;

architecture SYN_ARCHSTRUCT of iv_8146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8145 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8145;

architecture SYN_ARCHSTRUCT of iv_8145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8144 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8144;

architecture SYN_ARCHSTRUCT of iv_8144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8143 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8143;

architecture SYN_ARCHSTRUCT of iv_8143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8142 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8142;

architecture SYN_ARCHSTRUCT of iv_8142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8141 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8141;

architecture SYN_ARCHSTRUCT of iv_8141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8140 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8140;

architecture SYN_ARCHSTRUCT of iv_8140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8139 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8139;

architecture SYN_ARCHSTRUCT of iv_8139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8138 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8138;

architecture SYN_ARCHSTRUCT of iv_8138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8137 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8137;

architecture SYN_ARCHSTRUCT of iv_8137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8136 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8136;

architecture SYN_ARCHSTRUCT of iv_8136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8135 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8135;

architecture SYN_ARCHSTRUCT of iv_8135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8134 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8134;

architecture SYN_ARCHSTRUCT of iv_8134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8133 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8133;

architecture SYN_ARCHSTRUCT of iv_8133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8132 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8132;

architecture SYN_ARCHSTRUCT of iv_8132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8131 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8131;

architecture SYN_ARCHSTRUCT of iv_8131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8130 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8130;

architecture SYN_ARCHSTRUCT of iv_8130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8129 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8129;

architecture SYN_ARCHSTRUCT of iv_8129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_251 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_251;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_251 is

   component muxN1_N4_251
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_501
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_502
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1096, n_1097 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_502 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1096);
   RCA2 : RCA_N4_501 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1097);
   MUX : muxN1_N4_251 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_250 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_250;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_250 is

   component muxN1_N4_250
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_499
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_500
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1098, n_1099 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_500 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1098);
   RCA2 : RCA_N4_499 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1099);
   MUX : muxN1_N4_250 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_249 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_249;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_249 is

   component muxN1_N4_249
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_497
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_498
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1100, n_1101 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_498 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1100);
   RCA2 : RCA_N4_497 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1101);
   MUX : muxN1_N4_249 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_248 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_248;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_248 is

   component muxN1_N4_248
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_495
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_496
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1102, n_1103 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_496 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1102);
   RCA2 : RCA_N4_495 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1103);
   MUX : muxN1_N4_248 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_247 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_247;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_247 is

   component muxN1_N4_247
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_493
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_494
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1104, n_1105 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_494 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1104);
   RCA2 : RCA_N4_493 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1105);
   MUX : muxN1_N4_247 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_246 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_246;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_246 is

   component muxN1_N4_246
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_491
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_492
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1106, n_1107 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_492 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1106);
   RCA2 : RCA_N4_491 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1107);
   MUX : muxN1_N4_246 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_245 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_245;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_245 is

   component muxN1_N4_245
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_489
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_490
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1108, n_1109 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_490 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1108);
   RCA2 : RCA_N4_489 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1109);
   MUX : muxN1_N4_245 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_244 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_244;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_244 is

   component muxN1_N4_244
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_487
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_488
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1110, n_1111 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_488 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1110);
   RCA2 : RCA_N4_487 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1111);
   MUX : muxN1_N4_244 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_243 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_243;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_243 is

   component muxN1_N4_243
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_485
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_486
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1112, n_1113 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_486 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1112);
   RCA2 : RCA_N4_485 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1113);
   MUX : muxN1_N4_243 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_242 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_242;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_242 is

   component muxN1_N4_242
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_483
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_484
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1114, n_1115 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_484 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1114);
   RCA2 : RCA_N4_483 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1115);
   MUX : muxN1_N4_242 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_241 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_241;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_241 is

   component muxN1_N4_241
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_481
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_482
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1116, n_1117 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_482 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1116);
   RCA2 : RCA_N4_481 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1117);
   MUX : muxN1_N4_241 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_generator_sparse_tree_N16_carry_range4_2 is

   port( P, G : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C : 
         out std_logic_vector (4 downto 0));

end carry_generator_sparse_tree_N16_carry_range4_2;

architecture SYN_ARCHSTRUCT of carry_generator_sparse_tree_N16_carry_range4_2 
   is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component g_block_261
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component g_block_262
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_957
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_263
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_958
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_959
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_960
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_264
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_961
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_962
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_963
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_964
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_965
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_966
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_967
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_265
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   signal C_4_port, C_3_port, C_2_port, C_1_port, Gmat_16_15_port, 
      Gmat_16_13_port, Gmat_16_9_port, Gmat_14_13_port, Gmat_12_11_port, 
      Gmat_12_9_port, Gmat_10_9_port, Gmat_8_7_port, Gmat_8_5_port, 
      Gmat_6_5_port, Gmat_4_3_port, Gmat_2_1_port, Pmat_16_15_port, 
      Pmat_16_13_port, Pmat_16_9_port, Pmat_14_13_port, Pmat_12_11_port, 
      Pmat_12_9_port, Pmat_10_9_port, Pmat_8_7_port, Pmat_8_5_port, 
      Pmat_6_5_port, Pmat_4_3_port, n1, n2 : std_logic;

begin
   C <= ( C_4_port, C_3_port, C_2_port, C_1_port, Cin );
   
   first_G_1_2 : g_block_265 port map( G_i_k => G(1), G_kmin1_j => n2, P_i_k =>
                           P(1), G_i_j => Gmat_2_1_port);
   FRST_PG_1_4 : pg_block_967 port map( G_i_k => G(3), G_kmin1_j => G(2), P_i_k
                           => P(3), P_kmin1_j => P(2), P_i_j => Pmat_4_3_port, 
                           G_i_j => Gmat_4_3_port);
   FRST_PG_1_6 : pg_block_966 port map( G_i_k => G(5), G_kmin1_j => G(4), P_i_k
                           => P(5), P_kmin1_j => P(4), P_i_j => Pmat_6_5_port, 
                           G_i_j => Gmat_6_5_port);
   FRST_PG_1_8 : pg_block_965 port map( G_i_k => G(7), G_kmin1_j => G(6), P_i_k
                           => P(7), P_kmin1_j => P(6), P_i_j => Pmat_8_7_port, 
                           G_i_j => Gmat_8_7_port);
   FRST_PG_1_10 : pg_block_964 port map( G_i_k => G(9), G_kmin1_j => G(8), 
                           P_i_k => P(9), P_kmin1_j => P(8), P_i_j => 
                           Pmat_10_9_port, G_i_j => Gmat_10_9_port);
   FRST_PG_1_12 : pg_block_963 port map( G_i_k => G(11), G_kmin1_j => G(10), 
                           P_i_k => P(11), P_kmin1_j => P(10), P_i_j => 
                           Pmat_12_11_port, G_i_j => Gmat_12_11_port);
   FRST_PG_1_14 : pg_block_962 port map( G_i_k => G(13), G_kmin1_j => G(12), 
                           P_i_k => P(13), P_kmin1_j => P(12), P_i_j => 
                           Pmat_14_13_port, G_i_j => Gmat_14_13_port);
   FRST_PG_1_16 : pg_block_961 port map( G_i_k => G(15), G_kmin1_j => G(14), 
                           P_i_k => P(15), P_kmin1_j => P(14), P_i_j => 
                           Pmat_16_15_port, G_i_j => Gmat_16_15_port);
   first_G_2_4 : g_block_264 port map( G_i_k => Gmat_4_3_port, G_kmin1_j => 
                           Gmat_2_1_port, P_i_k => Pmat_4_3_port, G_i_j => 
                           C_1_port);
   FRST_PG_2_8 : pg_block_960 port map( G_i_k => Gmat_8_7_port, G_kmin1_j => 
                           Gmat_6_5_port, P_i_k => Pmat_8_7_port, P_kmin1_j => 
                           Pmat_6_5_port, P_i_j => Pmat_8_5_port, G_i_j => 
                           Gmat_8_5_port);
   FRST_PG_2_12 : pg_block_959 port map( G_i_k => Gmat_12_11_port, G_kmin1_j =>
                           Gmat_10_9_port, P_i_k => Pmat_12_11_port, P_kmin1_j 
                           => Pmat_10_9_port, P_i_j => Pmat_12_9_port, G_i_j =>
                           Gmat_12_9_port);
   FRST_PG_2_16 : pg_block_958 port map( G_i_k => Gmat_16_15_port, G_kmin1_j =>
                           Gmat_14_13_port, P_i_k => Pmat_16_15_port, P_kmin1_j
                           => Pmat_14_13_port, P_i_j => Pmat_16_13_port, G_i_j 
                           => Gmat_16_13_port);
   G_L2_0_4_8 : g_block_263 port map( G_i_k => Gmat_8_5_port, G_kmin1_j => 
                           C_1_port, P_i_k => Pmat_8_5_port, G_i_j => C_2_port)
                           ;
   PG_L2_0_12_16 : pg_block_957 port map( G_i_k => Gmat_16_13_port, G_kmin1_j 
                           => Gmat_12_9_port, P_i_k => Pmat_16_13_port, 
                           P_kmin1_j => Pmat_12_9_port, P_i_j => Pmat_16_9_port
                           , G_i_j => Gmat_16_9_port);
   G_L2_1_8_12 : g_block_262 port map( G_i_k => Gmat_12_9_port, G_kmin1_j => 
                           C_2_port, P_i_k => Pmat_12_9_port, G_i_j => C_3_port
                           );
   G_L2_1_8_16 : g_block_261 port map( G_i_k => Gmat_16_9_port, G_kmin1_j => 
                           C_2_port, P_i_k => Pmat_16_9_port, G_i_j => C_4_port
                           );
   U1 : INV_X1 port map( A => n1, ZN => n2);
   U2 : AOI21_X1 port map( B1 => P(0), B2 => Cin, A => G(0), ZN => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_generator_sparse_tree_N16_carry_range4_1 is

   port( P, G : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C : 
         out std_logic_vector (4 downto 0));

end carry_generator_sparse_tree_N16_carry_range4_1;

architecture SYN_ARCHSTRUCT of carry_generator_sparse_tree_N16_carry_range4_1 
   is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component g_block_256
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component g_block_257
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_946
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_258
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_947
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_948
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_949
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_259
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_950
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_951
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_952
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_953
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_954
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_955
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_956
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_260
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   signal C_4_port, C_3_port, C_2_port, C_1_port, Gmat_16_15_port, 
      Gmat_16_13_port, Gmat_16_9_port, Gmat_14_13_port, Gmat_12_11_port, 
      Gmat_12_9_port, Gmat_10_9_port, Gmat_8_7_port, Gmat_8_5_port, 
      Gmat_6_5_port, Gmat_4_3_port, Gmat_2_1_port, Pmat_16_15_port, 
      Pmat_16_13_port, Pmat_16_9_port, Pmat_14_13_port, Pmat_12_11_port, 
      Pmat_12_9_port, Pmat_10_9_port, Pmat_8_7_port, Pmat_8_5_port, 
      Pmat_6_5_port, Pmat_4_3_port, n1, n2 : std_logic;

begin
   C <= ( C_4_port, C_3_port, C_2_port, C_1_port, Cin );
   
   first_G_1_2 : g_block_260 port map( G_i_k => G(1), G_kmin1_j => n2, P_i_k =>
                           P(1), G_i_j => Gmat_2_1_port);
   FRST_PG_1_4 : pg_block_956 port map( G_i_k => G(3), G_kmin1_j => G(2), P_i_k
                           => P(3), P_kmin1_j => P(2), P_i_j => Pmat_4_3_port, 
                           G_i_j => Gmat_4_3_port);
   FRST_PG_1_6 : pg_block_955 port map( G_i_k => G(5), G_kmin1_j => G(4), P_i_k
                           => P(5), P_kmin1_j => P(4), P_i_j => Pmat_6_5_port, 
                           G_i_j => Gmat_6_5_port);
   FRST_PG_1_8 : pg_block_954 port map( G_i_k => G(7), G_kmin1_j => G(6), P_i_k
                           => P(7), P_kmin1_j => P(6), P_i_j => Pmat_8_7_port, 
                           G_i_j => Gmat_8_7_port);
   FRST_PG_1_10 : pg_block_953 port map( G_i_k => G(9), G_kmin1_j => G(8), 
                           P_i_k => P(9), P_kmin1_j => P(8), P_i_j => 
                           Pmat_10_9_port, G_i_j => Gmat_10_9_port);
   FRST_PG_1_12 : pg_block_952 port map( G_i_k => G(11), G_kmin1_j => G(10), 
                           P_i_k => P(11), P_kmin1_j => P(10), P_i_j => 
                           Pmat_12_11_port, G_i_j => Gmat_12_11_port);
   FRST_PG_1_14 : pg_block_951 port map( G_i_k => G(13), G_kmin1_j => G(12), 
                           P_i_k => P(13), P_kmin1_j => P(12), P_i_j => 
                           Pmat_14_13_port, G_i_j => Gmat_14_13_port);
   FRST_PG_1_16 : pg_block_950 port map( G_i_k => G(15), G_kmin1_j => G(14), 
                           P_i_k => P(15), P_kmin1_j => P(14), P_i_j => 
                           Pmat_16_15_port, G_i_j => Gmat_16_15_port);
   first_G_2_4 : g_block_259 port map( G_i_k => Gmat_4_3_port, G_kmin1_j => 
                           Gmat_2_1_port, P_i_k => Pmat_4_3_port, G_i_j => 
                           C_1_port);
   FRST_PG_2_8 : pg_block_949 port map( G_i_k => Gmat_8_7_port, G_kmin1_j => 
                           Gmat_6_5_port, P_i_k => Pmat_8_7_port, P_kmin1_j => 
                           Pmat_6_5_port, P_i_j => Pmat_8_5_port, G_i_j => 
                           Gmat_8_5_port);
   FRST_PG_2_12 : pg_block_948 port map( G_i_k => Gmat_12_11_port, G_kmin1_j =>
                           Gmat_10_9_port, P_i_k => Pmat_12_11_port, P_kmin1_j 
                           => Pmat_10_9_port, P_i_j => Pmat_12_9_port, G_i_j =>
                           Gmat_12_9_port);
   FRST_PG_2_16 : pg_block_947 port map( G_i_k => Gmat_16_15_port, G_kmin1_j =>
                           Gmat_14_13_port, P_i_k => Pmat_16_15_port, P_kmin1_j
                           => Pmat_14_13_port, P_i_j => Pmat_16_13_port, G_i_j 
                           => Gmat_16_13_port);
   G_L2_0_4_8 : g_block_258 port map( G_i_k => Gmat_8_5_port, G_kmin1_j => 
                           C_1_port, P_i_k => Pmat_8_5_port, G_i_j => C_2_port)
                           ;
   PG_L2_0_12_16 : pg_block_946 port map( G_i_k => Gmat_16_13_port, G_kmin1_j 
                           => Gmat_12_9_port, P_i_k => Pmat_16_13_port, 
                           P_kmin1_j => Pmat_12_9_port, P_i_j => Pmat_16_9_port
                           , G_i_j => Gmat_16_9_port);
   G_L2_1_8_12 : g_block_257 port map( G_i_k => Gmat_12_9_port, G_kmin1_j => 
                           C_2_port, P_i_k => Pmat_12_9_port, G_i_j => C_3_port
                           );
   G_L2_1_8_16 : g_block_256 port map( G_i_k => Gmat_16_9_port, G_kmin1_j => 
                           C_2_port, P_i_k => Pmat_16_9_port, G_i_j => C_4_port
                           );
   U1 : INV_X1 port map( A => n1, ZN => n2);
   U2 : AOI21_X1 port map( B1 => P(0), B2 => Cin, A => G(0), ZN => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_network_N16_2 is

   port( A, B : in std_logic_vector (15 downto 0);  P, G : out std_logic_vector
         (15 downto 0));

end pg_network_N16_2;

architecture SYN_ARCHDATAFLOW of pg_network_N16_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B(9), B => A(9), Z => P(9));
   U2 : XOR2_X1 port map( A => B(8), B => A(8), Z => P(8));
   U3 : XOR2_X1 port map( A => B(7), B => A(7), Z => P(7));
   U4 : XOR2_X1 port map( A => B(6), B => A(6), Z => P(6));
   U5 : XOR2_X1 port map( A => B(5), B => A(5), Z => P(5));
   U6 : XOR2_X1 port map( A => B(4), B => A(4), Z => P(4));
   U7 : XOR2_X1 port map( A => B(3), B => A(3), Z => P(3));
   U8 : XOR2_X1 port map( A => B(2), B => A(2), Z => P(2));
   U9 : XOR2_X1 port map( A => B(1), B => A(1), Z => P(1));
   U10 : XOR2_X1 port map( A => B(15), B => A(15), Z => P(15));
   U11 : XOR2_X1 port map( A => B(14), B => A(14), Z => P(14));
   U12 : XOR2_X1 port map( A => B(13), B => A(13), Z => P(13));
   U13 : XOR2_X1 port map( A => B(12), B => A(12), Z => P(12));
   U14 : XOR2_X1 port map( A => B(11), B => A(11), Z => P(11));
   U15 : XOR2_X1 port map( A => B(10), B => A(10), Z => P(10));
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => P(0));
   U17 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => G(9));
   U18 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => G(8));
   U19 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => G(7));
   U20 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => G(6));
   U21 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => G(5));
   U22 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => G(4));
   U23 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => G(3));
   U24 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => G(2));
   U25 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => G(1));
   U26 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => G(15));
   U27 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => G(14));
   U28 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => G(13));
   U29 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => G(12));
   U30 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => G(11));
   U31 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => G(10));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => G(0));

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_network_N16_1 is

   port( A, B : in std_logic_vector (15 downto 0);  P, G : out std_logic_vector
         (15 downto 0));

end pg_network_N16_1;

architecture SYN_ARCHDATAFLOW of pg_network_N16_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B(9), B => A(9), Z => P(9));
   U2 : XOR2_X1 port map( A => B(8), B => A(8), Z => P(8));
   U3 : XOR2_X1 port map( A => B(7), B => A(7), Z => P(7));
   U4 : XOR2_X1 port map( A => B(6), B => A(6), Z => P(6));
   U5 : XOR2_X1 port map( A => B(5), B => A(5), Z => P(5));
   U6 : XOR2_X1 port map( A => B(4), B => A(4), Z => P(4));
   U7 : XOR2_X1 port map( A => B(3), B => A(3), Z => P(3));
   U8 : XOR2_X1 port map( A => B(2), B => A(2), Z => P(2));
   U9 : XOR2_X1 port map( A => B(1), B => A(1), Z => P(1));
   U10 : XOR2_X1 port map( A => B(15), B => A(15), Z => P(15));
   U11 : XOR2_X1 port map( A => B(14), B => A(14), Z => P(14));
   U12 : XOR2_X1 port map( A => B(13), B => A(13), Z => P(13));
   U13 : XOR2_X1 port map( A => B(12), B => A(12), Z => P(12));
   U14 : XOR2_X1 port map( A => B(11), B => A(11), Z => P(11));
   U15 : XOR2_X1 port map( A => B(10), B => A(10), Z => P(10));
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => P(0));
   U17 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => G(9));
   U18 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => G(8));
   U19 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => G(7));
   U20 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => G(6));
   U21 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => G(5));
   U22 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => G(4));
   U23 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => G(3));
   U24 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => G(2));
   U25 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => G(1));
   U26 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => G(15));
   U27 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => G(14));
   U28 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => G(13));
   U29 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => G(12));
   U30 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => G(11));
   U31 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => G(10));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => G(0));

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8623 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8623;

architecture SYN_ARCHSTRUCT of mux21_8623 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25867
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25868
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25869
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8623
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8623 port map( A => n1, Y => n_S);
   NAND1 : nd2_25869 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25868 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25867 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8622 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8622;

architecture SYN_ARCHSTRUCT of mux21_8622 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25864
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25865
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25866
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8622
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8622 port map( A => n1, Y => n_S);
   NAND1 : nd2_25866 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25865 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25864 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8621 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8621;

architecture SYN_ARCHSTRUCT of mux21_8621 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25861
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25862
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25863
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8621
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8621 port map( A => n1, Y => n_S);
   NAND1 : nd2_25863 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25862 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25861 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8620 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8620;

architecture SYN_ARCHSTRUCT of mux21_8620 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25858
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25859
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25860
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8620
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8620 port map( A => n1, Y => n_S);
   NAND1 : nd2_25860 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25859 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25858 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8619 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8619;

architecture SYN_ARCHSTRUCT of mux21_8619 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25855
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25856
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25857
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8619
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8619 port map( A => n1, Y => n_S);
   NAND1 : nd2_25857 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25856 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25855 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8618 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8618;

architecture SYN_ARCHSTRUCT of mux21_8618 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25852
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25853
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25854
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8618
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8618 port map( A => n1, Y => n_S);
   NAND1 : nd2_25854 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25853 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25852 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8617 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8617;

architecture SYN_ARCHSTRUCT of mux21_8617 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25849
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25850
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25851
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8617
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8617 port map( A => n1, Y => n_S);
   NAND1 : nd2_25851 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25850 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25849 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8616 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8616;

architecture SYN_ARCHSTRUCT of mux21_8616 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25846
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25847
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25848
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8616
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8616 port map( A => n1, Y => n_S);
   NAND1 : nd2_25848 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25847 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25846 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8615 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8615;

architecture SYN_ARCHSTRUCT of mux21_8615 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25843
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25844
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25845
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8615
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8615 port map( A => n1, Y => n_S);
   NAND1 : nd2_25845 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25844 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25843 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8614 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8614;

architecture SYN_ARCHSTRUCT of mux21_8614 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25840
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25841
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25842
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8614
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8614 port map( A => n1, Y => n_S);
   NAND1 : nd2_25842 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25841 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25840 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8613 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8613;

architecture SYN_ARCHSTRUCT of mux21_8613 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25837
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25838
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25839
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8613
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8613 port map( A => n1, Y => n_S);
   NAND1 : nd2_25839 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25838 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25837 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8612 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8612;

architecture SYN_ARCHSTRUCT of mux21_8612 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25834
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25835
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25836
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8612
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8612 port map( A => n1, Y => n_S);
   NAND1 : nd2_25836 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25835 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25834 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8611 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8611;

architecture SYN_ARCHSTRUCT of mux21_8611 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25831
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25832
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25833
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8611
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8611 port map( A => n1, Y => n_S);
   NAND1 : nd2_25833 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25832 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25831 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8610 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8610;

architecture SYN_ARCHSTRUCT of mux21_8610 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25828
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25829
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25830
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8610
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8610 port map( A => n1, Y => n_S);
   NAND1 : nd2_25830 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25829 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25828 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8609 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8609;

architecture SYN_ARCHSTRUCT of mux21_8609 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25825
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25826
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25827
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8609
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8609 port map( A => n1, Y => n_S);
   NAND1 : nd2_25827 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25826 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25825 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8608 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8608;

architecture SYN_ARCHSTRUCT of mux21_8608 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25822
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25823
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25824
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8608
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8608 port map( A => n1, Y => n_S);
   NAND1 : nd2_25824 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25823 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25822 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8607 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8607;

architecture SYN_ARCHSTRUCT of mux21_8607 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25819
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25820
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25821
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8607
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8607 port map( A => n1, Y => n_S);
   NAND1 : nd2_25821 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25820 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25819 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8606 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8606;

architecture SYN_ARCHSTRUCT of mux21_8606 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25816
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25817
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25818
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8606
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8606 port map( A => n1, Y => n_S);
   NAND1 : nd2_25818 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25817 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25816 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8605 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8605;

architecture SYN_ARCHSTRUCT of mux21_8605 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25813
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25814
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25815
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8605
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8605 port map( A => n1, Y => n_S);
   NAND1 : nd2_25815 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25814 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25813 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8604 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8604;

architecture SYN_ARCHSTRUCT of mux21_8604 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25810
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25811
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25812
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8604
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8604 port map( A => n1, Y => n_S);
   NAND1 : nd2_25812 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25811 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25810 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8603 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8603;

architecture SYN_ARCHSTRUCT of mux21_8603 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25807
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25808
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25809
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8603
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8603 port map( A => n1, Y => n_S);
   NAND1 : nd2_25809 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25808 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25807 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8602 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8602;

architecture SYN_ARCHSTRUCT of mux21_8602 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25804
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25805
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25806
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8602
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8602 port map( A => n1, Y => n_S);
   NAND1 : nd2_25806 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25805 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25804 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8601 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8601;

architecture SYN_ARCHSTRUCT of mux21_8601 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25801
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25802
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25803
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8601
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8601 port map( A => n1, Y => n_S);
   NAND1 : nd2_25803 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25802 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25801 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8600 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8600;

architecture SYN_ARCHSTRUCT of mux21_8600 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25798
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25799
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25800
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8600
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8600 port map( A => n1, Y => n_S);
   NAND1 : nd2_25800 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25799 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25798 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8599 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8599;

architecture SYN_ARCHSTRUCT of mux21_8599 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25795
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25796
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25797
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8599
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8599 port map( A => n1, Y => n_S);
   NAND1 : nd2_25797 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25796 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25795 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8598 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8598;

architecture SYN_ARCHSTRUCT of mux21_8598 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25792
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25793
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25794
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8598
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8598 port map( A => n1, Y => n_S);
   NAND1 : nd2_25794 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25793 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25792 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8597 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8597;

architecture SYN_ARCHSTRUCT of mux21_8597 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25789
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25790
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25791
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8597
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8597 port map( A => n1, Y => n_S);
   NAND1 : nd2_25791 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25790 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25789 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8596 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8596;

architecture SYN_ARCHSTRUCT of mux21_8596 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25786
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25787
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25788
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8596
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8596 port map( A => n1, Y => n_S);
   NAND1 : nd2_25788 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25787 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25786 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8595 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8595;

architecture SYN_ARCHSTRUCT of mux21_8595 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25783
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25784
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25785
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8595
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8595 port map( A => n1, Y => n_S);
   NAND1 : nd2_25785 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25784 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25783 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8594 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8594;

architecture SYN_ARCHSTRUCT of mux21_8594 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25780
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25781
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25782
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8594
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8594 port map( A => n1, Y => n_S);
   NAND1 : nd2_25782 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25781 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25780 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8593 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8593;

architecture SYN_ARCHSTRUCT of mux21_8593 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25777
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25778
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25779
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8593
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8593 port map( A => n1, Y => n_S);
   NAND1 : nd2_25779 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25778 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25777 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8592 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8592;

architecture SYN_ARCHSTRUCT of mux21_8592 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25774
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25775
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25776
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8592
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8592 port map( A => n1, Y => n_S);
   NAND1 : nd2_25776 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25775 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25774 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8591 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8591;

architecture SYN_ARCHSTRUCT of mux21_8591 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25771
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25772
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25773
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8591
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8591 port map( A => n1, Y => n_S);
   NAND1 : nd2_25773 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25772 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25771 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8590 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8590;

architecture SYN_ARCHSTRUCT of mux21_8590 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25768
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25769
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25770
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8590
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8590 port map( A => n1, Y => n_S);
   NAND1 : nd2_25770 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25769 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25768 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8589 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8589;

architecture SYN_ARCHSTRUCT of mux21_8589 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25765
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25766
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25767
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8589
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8589 port map( A => n1, Y => n_S);
   NAND1 : nd2_25767 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25766 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25765 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8588 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8588;

architecture SYN_ARCHSTRUCT of mux21_8588 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25762
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25763
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25764
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8588
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8588 port map( A => n1, Y => n_S);
   NAND1 : nd2_25764 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25763 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25762 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8587 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8587;

architecture SYN_ARCHSTRUCT of mux21_8587 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25759
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25760
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25761
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8587
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8587 port map( A => n1, Y => n_S);
   NAND1 : nd2_25761 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25760 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25759 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8586 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8586;

architecture SYN_ARCHSTRUCT of mux21_8586 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25756
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25757
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25758
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8586
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8586 port map( A => n1, Y => n_S);
   NAND1 : nd2_25758 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25757 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25756 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8585 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8585;

architecture SYN_ARCHSTRUCT of mux21_8585 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25753
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25754
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25755
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8585
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8585 port map( A => n1, Y => n_S);
   NAND1 : nd2_25755 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25754 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25753 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8584 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8584;

architecture SYN_ARCHSTRUCT of mux21_8584 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25750
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25751
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25752
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8584
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8584 port map( A => n1, Y => n_S);
   NAND1 : nd2_25752 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25751 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25750 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8583 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8583;

architecture SYN_ARCHSTRUCT of mux21_8583 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25747
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25748
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25749
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8583
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8583 port map( A => n1, Y => n_S);
   NAND1 : nd2_25749 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25748 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25747 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8582 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8582;

architecture SYN_ARCHSTRUCT of mux21_8582 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25744
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25745
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25746
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8582
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8582 port map( A => n1, Y => n_S);
   NAND1 : nd2_25746 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25745 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25744 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8581 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8581;

architecture SYN_ARCHSTRUCT of mux21_8581 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25741
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25742
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25743
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8581
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8581 port map( A => n1, Y => n_S);
   NAND1 : nd2_25743 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25742 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25741 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8580 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8580;

architecture SYN_ARCHSTRUCT of mux21_8580 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25738
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25739
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25740
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8580
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8580 port map( A => n1, Y => n_S);
   NAND1 : nd2_25740 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25739 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25738 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8579 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8579;

architecture SYN_ARCHSTRUCT of mux21_8579 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25735
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25736
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25737
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8579
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8579 port map( A => n1, Y => n_S);
   NAND1 : nd2_25737 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25736 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25735 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8578 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8578;

architecture SYN_ARCHSTRUCT of mux21_8578 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25732
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25733
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25734
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8578
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8578 port map( A => n1, Y => n_S);
   NAND1 : nd2_25734 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25733 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25732 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8577 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8577;

architecture SYN_ARCHSTRUCT of mux21_8577 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25729
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25730
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25731
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8577
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8577 port map( A => n1, Y => n_S);
   NAND1 : nd2_25731 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25730 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25729 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8576 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8576;

architecture SYN_ARCHSTRUCT of mux21_8576 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25726
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25727
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25728
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8576
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8576 port map( A => n1, Y => n_S);
   NAND1 : nd2_25728 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25727 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25726 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8575 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8575;

architecture SYN_ARCHSTRUCT of mux21_8575 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25723
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25724
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25725
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8575
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8575 port map( A => n1, Y => n_S);
   NAND1 : nd2_25725 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25724 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25723 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8574 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8574;

architecture SYN_ARCHSTRUCT of mux21_8574 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25720
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25721
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25722
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8574
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8574 port map( A => n1, Y => n_S);
   NAND1 : nd2_25722 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25721 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25720 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8573 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8573;

architecture SYN_ARCHSTRUCT of mux21_8573 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25717
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25718
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25719
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8573
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8573 port map( A => n1, Y => n_S);
   NAND1 : nd2_25719 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25718 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25717 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8572 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8572;

architecture SYN_ARCHSTRUCT of mux21_8572 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25714
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25715
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25716
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8572
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8572 port map( A => n1, Y => n_S);
   NAND1 : nd2_25716 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25715 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25714 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8571 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8571;

architecture SYN_ARCHSTRUCT of mux21_8571 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25711
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25712
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25713
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8571
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8571 port map( A => n1, Y => n_S);
   NAND1 : nd2_25713 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25712 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25711 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8570 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8570;

architecture SYN_ARCHSTRUCT of mux21_8570 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25708
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25709
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25710
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8570
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8570 port map( A => n1, Y => n_S);
   NAND1 : nd2_25710 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25709 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25708 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8569 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8569;

architecture SYN_ARCHSTRUCT of mux21_8569 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25705
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25706
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25707
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8569
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8569 port map( A => n1, Y => n_S);
   NAND1 : nd2_25707 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25706 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25705 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8568 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8568;

architecture SYN_ARCHSTRUCT of mux21_8568 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25702
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25703
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25704
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8568
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8568 port map( A => n1, Y => n_S);
   NAND1 : nd2_25704 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25703 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25702 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8567 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8567;

architecture SYN_ARCHSTRUCT of mux21_8567 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25699
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25700
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25701
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8567
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8567 port map( A => n1, Y => n_S);
   NAND1 : nd2_25701 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25700 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25699 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8566 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8566;

architecture SYN_ARCHSTRUCT of mux21_8566 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25696
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25697
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25698
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8566
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8566 port map( A => n1, Y => n_S);
   NAND1 : nd2_25698 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25697 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25696 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8565 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8565;

architecture SYN_ARCHSTRUCT of mux21_8565 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25693
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25694
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25695
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8565
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8565 port map( A => n1, Y => n_S);
   NAND1 : nd2_25695 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25694 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25693 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8564 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8564;

architecture SYN_ARCHSTRUCT of mux21_8564 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25690
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25691
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25692
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8564
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8564 port map( A => n1, Y => n_S);
   NAND1 : nd2_25692 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25691 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25690 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8563 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8563;

architecture SYN_ARCHSTRUCT of mux21_8563 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25687
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25688
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25689
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8563
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8563 port map( A => n1, Y => n_S);
   NAND1 : nd2_25689 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25688 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25687 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8562 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8562;

architecture SYN_ARCHSTRUCT of mux21_8562 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25684
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25685
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25686
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8562
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8562 port map( A => n1, Y => n_S);
   NAND1 : nd2_25686 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25685 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25684 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8561 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8561;

architecture SYN_ARCHSTRUCT of mux21_8561 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25681
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25682
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25683
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8561
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8561 port map( A => n1, Y => n_S);
   NAND1 : nd2_25683 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25682 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25681 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8560 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8560;

architecture SYN_ARCHSTRUCT of mux21_8560 is

   component nd2_25678
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25679
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25680
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8560
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8560 port map( A => S, Y => n_S);
   NAND1 : nd2_25680 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25679 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25678 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8559 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8559;

architecture SYN_ARCHSTRUCT of mux21_8559 is

   component nd2_25675
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25676
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25677
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8559
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8559 port map( A => S, Y => n_S);
   NAND1 : nd2_25677 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25676 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25675 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8558 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8558;

architecture SYN_ARCHSTRUCT of mux21_8558 is

   component nd2_25672
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25673
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25674
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8558
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8558 port map( A => S, Y => n_S);
   NAND1 : nd2_25674 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25673 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25672 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8557 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8557;

architecture SYN_ARCHSTRUCT of mux21_8557 is

   component nd2_25669
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25670
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25671
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8557
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8557 port map( A => S, Y => n_S);
   NAND1 : nd2_25671 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25670 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25669 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8556 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8556;

architecture SYN_ARCHSTRUCT of mux21_8556 is

   component nd2_25666
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25667
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25668
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8556
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8556 port map( A => S, Y => n_S);
   NAND1 : nd2_25668 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25667 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25666 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8555 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8555;

architecture SYN_ARCHSTRUCT of mux21_8555 is

   component nd2_25663
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25664
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25665
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8555
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8555 port map( A => S, Y => n_S);
   NAND1 : nd2_25665 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25664 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25663 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8554 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8554;

architecture SYN_ARCHSTRUCT of mux21_8554 is

   component nd2_25660
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25661
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25662
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8554
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8554 port map( A => S, Y => n_S);
   NAND1 : nd2_25662 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25661 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25660 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8553 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8553;

architecture SYN_ARCHSTRUCT of mux21_8553 is

   component nd2_25657
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25658
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25659
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8553
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8553 port map( A => S, Y => n_S);
   NAND1 : nd2_25659 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25658 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25657 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8552 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8552;

architecture SYN_ARCHSTRUCT of mux21_8552 is

   component nd2_25654
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25655
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25656
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8552
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8552 port map( A => S, Y => n_S);
   NAND1 : nd2_25656 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25655 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25654 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8551 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8551;

architecture SYN_ARCHSTRUCT of mux21_8551 is

   component nd2_25651
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25652
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25653
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8551
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8551 port map( A => S, Y => n_S);
   NAND1 : nd2_25653 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25652 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25651 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8550 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8550;

architecture SYN_ARCHSTRUCT of mux21_8550 is

   component nd2_25648
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25649
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25650
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8550
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8550 port map( A => S, Y => n_S);
   NAND1 : nd2_25650 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25649 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25648 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8549 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8549;

architecture SYN_ARCHSTRUCT of mux21_8549 is

   component nd2_25645
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25646
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25647
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8549
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8549 port map( A => S, Y => n_S);
   NAND1 : nd2_25647 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25646 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25645 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8548 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8548;

architecture SYN_ARCHSTRUCT of mux21_8548 is

   component nd2_25642
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25643
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25644
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8548
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8548 port map( A => S, Y => n_S);
   NAND1 : nd2_25644 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25643 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25642 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8547 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8547;

architecture SYN_ARCHSTRUCT of mux21_8547 is

   component nd2_25639
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25640
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25641
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8547
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8547 port map( A => S, Y => n_S);
   NAND1 : nd2_25641 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25640 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25639 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8546 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8546;

architecture SYN_ARCHSTRUCT of mux21_8546 is

   component nd2_25636
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25637
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25638
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8546
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8546 port map( A => S, Y => n_S);
   NAND1 : nd2_25638 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25637 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25636 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8545 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8545;

architecture SYN_ARCHSTRUCT of mux21_8545 is

   component nd2_25633
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25634
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25635
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8545
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8545 port map( A => S, Y => n_S);
   NAND1 : nd2_25635 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25634 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25633 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8544 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8544;

architecture SYN_ARCHSTRUCT of mux21_8544 is

   component nd2_25630
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25631
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25632
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8544
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8544 port map( A => S, Y => n_S);
   NAND1 : nd2_25632 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25631 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25630 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8543 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8543;

architecture SYN_ARCHSTRUCT of mux21_8543 is

   component nd2_25627
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25628
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25629
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8543
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8543 port map( A => S, Y => n_S);
   NAND1 : nd2_25629 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25628 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25627 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8542 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8542;

architecture SYN_ARCHSTRUCT of mux21_8542 is

   component nd2_25624
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25625
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25626
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8542
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8542 port map( A => S, Y => n_S);
   NAND1 : nd2_25626 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25625 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25624 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8541 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8541;

architecture SYN_ARCHSTRUCT of mux21_8541 is

   component nd2_25621
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25622
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25623
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8541
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8541 port map( A => S, Y => n_S);
   NAND1 : nd2_25623 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25622 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25621 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8540 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8540;

architecture SYN_ARCHSTRUCT of mux21_8540 is

   component nd2_25618
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25619
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25620
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8540
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8540 port map( A => S, Y => n_S);
   NAND1 : nd2_25620 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25619 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25618 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8539 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8539;

architecture SYN_ARCHSTRUCT of mux21_8539 is

   component nd2_25615
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25616
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25617
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8539
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8539 port map( A => S, Y => n_S);
   NAND1 : nd2_25617 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25616 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25615 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8538 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8538;

architecture SYN_ARCHSTRUCT of mux21_8538 is

   component nd2_25612
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25613
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25614
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8538
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8538 port map( A => S, Y => n_S);
   NAND1 : nd2_25614 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25613 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25612 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8537 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8537;

architecture SYN_ARCHSTRUCT of mux21_8537 is

   component nd2_25609
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25610
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25611
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8537
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8537 port map( A => S, Y => n_S);
   NAND1 : nd2_25611 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25610 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25609 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8536 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8536;

architecture SYN_ARCHSTRUCT of mux21_8536 is

   component nd2_25606
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25607
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25608
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8536
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8536 port map( A => S, Y => n_S);
   NAND1 : nd2_25608 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25607 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25606 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8535 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8535;

architecture SYN_ARCHSTRUCT of mux21_8535 is

   component nd2_25603
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25604
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25605
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8535
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8535 port map( A => S, Y => n_S);
   NAND1 : nd2_25605 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25604 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25603 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8534 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8534;

architecture SYN_ARCHSTRUCT of mux21_8534 is

   component nd2_25600
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25601
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25602
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8534
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8534 port map( A => S, Y => n_S);
   NAND1 : nd2_25602 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25601 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25600 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8533 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8533;

architecture SYN_ARCHSTRUCT of mux21_8533 is

   component nd2_25597
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25598
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25599
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8533
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8533 port map( A => S, Y => n_S);
   NAND1 : nd2_25599 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25598 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25597 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8532 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8532;

architecture SYN_ARCHSTRUCT of mux21_8532 is

   component nd2_25594
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25595
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25596
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8532
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8532 port map( A => S, Y => n_S);
   NAND1 : nd2_25596 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25595 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25594 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8531 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8531;

architecture SYN_ARCHSTRUCT of mux21_8531 is

   component nd2_25591
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25592
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25593
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8531
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8531 port map( A => S, Y => n_S);
   NAND1 : nd2_25593 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25592 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25591 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8530 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8530;

architecture SYN_ARCHSTRUCT of mux21_8530 is

   component nd2_25588
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25589
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25590
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8530
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8530 port map( A => S, Y => n_S);
   NAND1 : nd2_25590 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25589 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25588 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8529 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8529;

architecture SYN_ARCHSTRUCT of mux21_8529 is

   component nd2_25585
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25586
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25587
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8529
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8529 port map( A => S, Y => n_S);
   NAND1 : nd2_25587 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25586 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25585 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8528 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8528;

architecture SYN_ARCHSTRUCT of mux21_8528 is

   component nd2_25582
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25583
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25584
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8528
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8528 port map( A => S, Y => n_S);
   NAND1 : nd2_25584 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25583 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25582 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8527 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8527;

architecture SYN_ARCHSTRUCT of mux21_8527 is

   component nd2_25579
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25580
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25581
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8527
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8527 port map( A => S, Y => n_S);
   NAND1 : nd2_25581 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25580 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25579 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8526 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8526;

architecture SYN_ARCHSTRUCT of mux21_8526 is

   component nd2_25576
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25577
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25578
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8526
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8526 port map( A => S, Y => n_S);
   NAND1 : nd2_25578 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25577 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25576 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8525 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8525;

architecture SYN_ARCHSTRUCT of mux21_8525 is

   component nd2_25573
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25574
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25575
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8525
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8525 port map( A => S, Y => n_S);
   NAND1 : nd2_25575 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25574 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25573 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8524 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8524;

architecture SYN_ARCHSTRUCT of mux21_8524 is

   component nd2_25570
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25571
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25572
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8524
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8524 port map( A => S, Y => n_S);
   NAND1 : nd2_25572 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25571 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25570 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8523 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8523;

architecture SYN_ARCHSTRUCT of mux21_8523 is

   component nd2_25567
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25568
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25569
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8523
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8523 port map( A => S, Y => n_S);
   NAND1 : nd2_25569 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25568 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25567 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8522 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8522;

architecture SYN_ARCHSTRUCT of mux21_8522 is

   component nd2_25564
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25565
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25566
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8522
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8522 port map( A => S, Y => n_S);
   NAND1 : nd2_25566 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25565 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25564 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8521 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8521;

architecture SYN_ARCHSTRUCT of mux21_8521 is

   component nd2_25561
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25562
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25563
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8521
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8521 port map( A => S, Y => n_S);
   NAND1 : nd2_25563 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25562 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25561 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8520 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8520;

architecture SYN_ARCHSTRUCT of mux21_8520 is

   component nd2_25558
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25559
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25560
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8520
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8520 port map( A => S, Y => n_S);
   NAND1 : nd2_25560 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25559 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25558 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8519 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8519;

architecture SYN_ARCHSTRUCT of mux21_8519 is

   component nd2_25555
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25556
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25557
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8519
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8519 port map( A => S, Y => n_S);
   NAND1 : nd2_25557 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25556 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25555 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8518 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8518;

architecture SYN_ARCHSTRUCT of mux21_8518 is

   component nd2_25552
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25553
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25554
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8518
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8518 port map( A => S, Y => n_S);
   NAND1 : nd2_25554 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25553 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25552 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8517 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8517;

architecture SYN_ARCHSTRUCT of mux21_8517 is

   component nd2_25549
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25550
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25551
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8517
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8517 port map( A => S, Y => n_S);
   NAND1 : nd2_25551 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25550 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25549 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8516 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8516;

architecture SYN_ARCHSTRUCT of mux21_8516 is

   component nd2_25546
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25547
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25548
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8516
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8516 port map( A => S, Y => n_S);
   NAND1 : nd2_25548 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25547 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25546 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8515 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8515;

architecture SYN_ARCHSTRUCT of mux21_8515 is

   component nd2_25543
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25544
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25545
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8515
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8515 port map( A => S, Y => n_S);
   NAND1 : nd2_25545 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25544 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25543 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8514 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8514;

architecture SYN_ARCHSTRUCT of mux21_8514 is

   component nd2_25540
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25541
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25542
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8514
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8514 port map( A => S, Y => n_S);
   NAND1 : nd2_25542 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25541 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25540 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8513 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8513;

architecture SYN_ARCHSTRUCT of mux21_8513 is

   component nd2_25537
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25538
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25539
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8513
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8513 port map( A => S, Y => n_S);
   NAND1 : nd2_25539 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25538 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25537 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8512 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8512;

architecture SYN_ARCHSTRUCT of mux21_8512 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25534
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25535
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25536
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8512
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8512 port map( A => n1, Y => n_S);
   NAND1 : nd2_25536 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25535 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25534 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8511 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8511;

architecture SYN_ARCHSTRUCT of mux21_8511 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25531
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25532
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25533
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8511
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8511 port map( A => n1, Y => n_S);
   NAND1 : nd2_25533 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25532 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25531 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8510 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8510;

architecture SYN_ARCHSTRUCT of mux21_8510 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25528
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25529
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25530
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8510
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8510 port map( A => n1, Y => n_S);
   NAND1 : nd2_25530 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25529 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25528 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8509 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8509;

architecture SYN_ARCHSTRUCT of mux21_8509 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25525
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25526
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25527
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8509
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8509 port map( A => n1, Y => n_S);
   NAND1 : nd2_25527 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25526 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25525 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8508 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8508;

architecture SYN_ARCHSTRUCT of mux21_8508 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25522
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25523
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25524
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8508
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8508 port map( A => n1, Y => n_S);
   NAND1 : nd2_25524 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25523 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25522 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8507 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8507;

architecture SYN_ARCHSTRUCT of mux21_8507 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25519
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25520
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25521
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8507
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8507 port map( A => n1, Y => n_S);
   NAND1 : nd2_25521 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25520 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25519 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8506 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8506;

architecture SYN_ARCHSTRUCT of mux21_8506 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25516
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25517
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25518
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8506
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8506 port map( A => n1, Y => n_S);
   NAND1 : nd2_25518 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25517 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25516 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8505 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8505;

architecture SYN_ARCHSTRUCT of mux21_8505 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25513
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25514
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25515
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8505
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8505 port map( A => n1, Y => n_S);
   NAND1 : nd2_25515 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25514 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25513 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8504 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8504;

architecture SYN_ARCHSTRUCT of mux21_8504 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25510
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25511
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25512
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8504
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8504 port map( A => n1, Y => n_S);
   NAND1 : nd2_25512 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25511 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25510 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8503 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8503;

architecture SYN_ARCHSTRUCT of mux21_8503 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25507
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25508
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25509
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8503
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8503 port map( A => n1, Y => n_S);
   NAND1 : nd2_25509 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25508 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25507 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8502 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8502;

architecture SYN_ARCHSTRUCT of mux21_8502 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25504
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25505
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25506
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8502
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8502 port map( A => n1, Y => n_S);
   NAND1 : nd2_25506 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25505 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25504 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8501 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8501;

architecture SYN_ARCHSTRUCT of mux21_8501 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25501
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25502
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25503
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8501
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8501 port map( A => n1, Y => n_S);
   NAND1 : nd2_25503 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25502 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25501 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8500 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8500;

architecture SYN_ARCHSTRUCT of mux21_8500 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25498
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25499
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25500
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8500
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8500 port map( A => n1, Y => n_S);
   NAND1 : nd2_25500 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25499 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25498 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8499 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8499;

architecture SYN_ARCHSTRUCT of mux21_8499 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25495
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25496
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25497
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8499
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8499 port map( A => n1, Y => n_S);
   NAND1 : nd2_25497 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25496 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25495 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8498 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8498;

architecture SYN_ARCHSTRUCT of mux21_8498 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25492
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25493
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25494
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8498
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8498 port map( A => n1, Y => n_S);
   NAND1 : nd2_25494 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25493 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25492 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8497 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8497;

architecture SYN_ARCHSTRUCT of mux21_8497 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25489
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25490
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25491
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8497
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8497 port map( A => n1, Y => n_S);
   NAND1 : nd2_25491 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25490 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25489 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8496 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8496;

architecture SYN_ARCHSTRUCT of mux21_8496 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25486
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25487
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25488
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8496
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8496 port map( A => n1, Y => n_S);
   NAND1 : nd2_25488 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25487 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25486 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8495 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8495;

architecture SYN_ARCHSTRUCT of mux21_8495 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25483
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25484
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25485
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8495
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8495 port map( A => n1, Y => n_S);
   NAND1 : nd2_25485 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25484 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25483 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8494 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8494;

architecture SYN_ARCHSTRUCT of mux21_8494 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25480
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25481
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25482
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8494
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8494 port map( A => n1, Y => n_S);
   NAND1 : nd2_25482 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25481 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25480 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8493 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8493;

architecture SYN_ARCHSTRUCT of mux21_8493 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25477
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25478
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25479
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8493
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8493 port map( A => n1, Y => n_S);
   NAND1 : nd2_25479 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25478 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25477 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8492 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8492;

architecture SYN_ARCHSTRUCT of mux21_8492 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25474
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25475
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25476
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8492
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8492 port map( A => n1, Y => n_S);
   NAND1 : nd2_25476 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25475 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25474 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8491 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8491;

architecture SYN_ARCHSTRUCT of mux21_8491 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25471
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25472
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25473
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8491
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8491 port map( A => n1, Y => n_S);
   NAND1 : nd2_25473 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25472 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25471 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8490 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8490;

architecture SYN_ARCHSTRUCT of mux21_8490 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25468
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25469
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25470
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8490
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8490 port map( A => n1, Y => n_S);
   NAND1 : nd2_25470 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25469 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25468 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8489 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8489;

architecture SYN_ARCHSTRUCT of mux21_8489 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25465
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25466
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25467
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8489
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8489 port map( A => n1, Y => n_S);
   NAND1 : nd2_25467 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25466 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25465 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8488 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8488;

architecture SYN_ARCHSTRUCT of mux21_8488 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25462
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25463
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25464
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8488
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8488 port map( A => n1, Y => n_S);
   NAND1 : nd2_25464 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25463 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25462 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8487 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8487;

architecture SYN_ARCHSTRUCT of mux21_8487 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25459
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25460
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25461
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8487
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8487 port map( A => n1, Y => n_S);
   NAND1 : nd2_25461 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25460 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25459 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8486 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8486;

architecture SYN_ARCHSTRUCT of mux21_8486 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25456
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25457
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25458
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8486
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8486 port map( A => n1, Y => n_S);
   NAND1 : nd2_25458 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25457 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25456 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8485 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8485;

architecture SYN_ARCHSTRUCT of mux21_8485 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25453
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25454
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25455
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8485
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8485 port map( A => n1, Y => n_S);
   NAND1 : nd2_25455 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25454 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25453 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8484 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8484;

architecture SYN_ARCHSTRUCT of mux21_8484 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25450
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25451
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25452
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8484
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8484 port map( A => n1, Y => n_S);
   NAND1 : nd2_25452 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25451 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25450 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8483 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8483;

architecture SYN_ARCHSTRUCT of mux21_8483 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25447
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25448
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25449
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8483
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8483 port map( A => n1, Y => n_S);
   NAND1 : nd2_25449 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25448 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25447 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8482 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8482;

architecture SYN_ARCHSTRUCT of mux21_8482 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25444
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25445
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25446
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8482
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8482 port map( A => n1, Y => n_S);
   NAND1 : nd2_25446 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25445 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25444 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8481 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8481;

architecture SYN_ARCHSTRUCT of mux21_8481 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25441
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25442
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25443
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8481
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8481 port map( A => n1, Y => n_S);
   NAND1 : nd2_25443 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25442 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25441 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8480 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8480;

architecture SYN_ARCHSTRUCT of mux21_8480 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25438
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25439
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25440
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8480
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8480 port map( A => n1, Y => n_S);
   NAND1 : nd2_25440 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25439 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25438 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8479 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8479;

architecture SYN_ARCHSTRUCT of mux21_8479 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25435
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25436
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25437
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8479
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8479 port map( A => n1, Y => n_S);
   NAND1 : nd2_25437 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25436 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25435 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8478 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8478;

architecture SYN_ARCHSTRUCT of mux21_8478 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25432
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25433
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25434
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8478
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8478 port map( A => n1, Y => n_S);
   NAND1 : nd2_25434 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25433 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25432 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8477 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8477;

architecture SYN_ARCHSTRUCT of mux21_8477 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25429
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25430
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25431
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8477
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8477 port map( A => n1, Y => n_S);
   NAND1 : nd2_25431 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25430 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25429 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8476 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8476;

architecture SYN_ARCHSTRUCT of mux21_8476 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25426
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25427
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25428
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8476
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8476 port map( A => n1, Y => n_S);
   NAND1 : nd2_25428 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25427 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25426 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8475 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8475;

architecture SYN_ARCHSTRUCT of mux21_8475 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25423
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25424
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25425
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8475
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8475 port map( A => n1, Y => n_S);
   NAND1 : nd2_25425 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25424 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25423 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8474 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8474;

architecture SYN_ARCHSTRUCT of mux21_8474 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25420
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25421
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25422
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8474
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8474 port map( A => n1, Y => n_S);
   NAND1 : nd2_25422 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25421 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25420 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8473 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8473;

architecture SYN_ARCHSTRUCT of mux21_8473 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25417
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25418
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25419
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8473
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8473 port map( A => n1, Y => n_S);
   NAND1 : nd2_25419 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25418 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25417 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8472 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8472;

architecture SYN_ARCHSTRUCT of mux21_8472 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25414
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25415
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25416
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8472
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8472 port map( A => n1, Y => n_S);
   NAND1 : nd2_25416 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25415 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25414 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8471 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8471;

architecture SYN_ARCHSTRUCT of mux21_8471 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25411
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25412
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25413
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8471
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8471 port map( A => n1, Y => n_S);
   NAND1 : nd2_25413 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25412 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25411 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8470 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8470;

architecture SYN_ARCHSTRUCT of mux21_8470 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25408
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25409
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25410
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8470
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8470 port map( A => n1, Y => n_S);
   NAND1 : nd2_25410 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25409 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25408 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8469 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8469;

architecture SYN_ARCHSTRUCT of mux21_8469 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25405
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25406
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25407
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8469
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8469 port map( A => n1, Y => n_S);
   NAND1 : nd2_25407 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25406 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25405 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8468 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8468;

architecture SYN_ARCHSTRUCT of mux21_8468 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25402
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25403
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25404
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8468
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8468 port map( A => n1, Y => n_S);
   NAND1 : nd2_25404 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25403 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25402 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8467 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8467;

architecture SYN_ARCHSTRUCT of mux21_8467 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25399
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25400
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25401
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8467
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8467 port map( A => n1, Y => n_S);
   NAND1 : nd2_25401 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25400 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25399 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8466 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8466;

architecture SYN_ARCHSTRUCT of mux21_8466 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25396
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25397
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25398
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8466
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8466 port map( A => n1, Y => n_S);
   NAND1 : nd2_25398 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25397 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25396 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8465 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8465;

architecture SYN_ARCHSTRUCT of mux21_8465 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25393
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25394
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25395
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8465
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8465 port map( A => n1, Y => n_S);
   NAND1 : nd2_25395 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25394 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25393 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8464 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8464;

architecture SYN_ARCHSTRUCT of mux21_8464 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25390
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25391
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25392
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8464
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8464 port map( A => n1, Y => n_S);
   NAND1 : nd2_25392 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25391 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25390 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8463 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8463;

architecture SYN_ARCHSTRUCT of mux21_8463 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25387
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25388
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25389
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8463
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8463 port map( A => n1, Y => n_S);
   NAND1 : nd2_25389 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25388 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25387 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8462 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8462;

architecture SYN_ARCHSTRUCT of mux21_8462 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25384
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25385
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25386
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8462
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8462 port map( A => n1, Y => n_S);
   NAND1 : nd2_25386 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25385 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25384 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8461 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8461;

architecture SYN_ARCHSTRUCT of mux21_8461 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25381
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25382
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25383
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8461
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8461 port map( A => n1, Y => n_S);
   NAND1 : nd2_25383 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25382 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25381 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8460 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8460;

architecture SYN_ARCHSTRUCT of mux21_8460 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25378
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25379
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25380
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8460
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8460 port map( A => n1, Y => n_S);
   NAND1 : nd2_25380 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25379 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25378 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8459 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8459;

architecture SYN_ARCHSTRUCT of mux21_8459 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25375
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25376
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25377
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8459
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8459 port map( A => n1, Y => n_S);
   NAND1 : nd2_25377 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25376 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25375 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8458 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8458;

architecture SYN_ARCHSTRUCT of mux21_8458 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25372
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25373
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25374
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8458
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8458 port map( A => n1, Y => n_S);
   NAND1 : nd2_25374 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25373 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25372 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8457 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8457;

architecture SYN_ARCHSTRUCT of mux21_8457 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25369
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25370
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25371
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8457
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8457 port map( A => n1, Y => n_S);
   NAND1 : nd2_25371 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25370 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25369 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8456 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8456;

architecture SYN_ARCHSTRUCT of mux21_8456 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25366
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25367
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25368
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8456
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8456 port map( A => n1, Y => n_S);
   NAND1 : nd2_25368 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25367 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25366 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8455 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8455;

architecture SYN_ARCHSTRUCT of mux21_8455 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25363
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25364
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25365
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8455
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8455 port map( A => n1, Y => n_S);
   NAND1 : nd2_25365 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25364 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25363 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8454 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8454;

architecture SYN_ARCHSTRUCT of mux21_8454 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25360
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25361
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25362
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8454
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8454 port map( A => n1, Y => n_S);
   NAND1 : nd2_25362 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25361 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25360 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8453 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8453;

architecture SYN_ARCHSTRUCT of mux21_8453 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25357
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25358
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25359
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8453
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8453 port map( A => n1, Y => n_S);
   NAND1 : nd2_25359 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25358 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25357 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8452 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8452;

architecture SYN_ARCHSTRUCT of mux21_8452 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25354
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25355
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25356
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8452
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8452 port map( A => n1, Y => n_S);
   NAND1 : nd2_25356 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25355 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25354 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8451 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8451;

architecture SYN_ARCHSTRUCT of mux21_8451 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25351
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25352
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25353
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8451
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8451 port map( A => n1, Y => n_S);
   NAND1 : nd2_25353 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25352 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25351 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8450 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8450;

architecture SYN_ARCHSTRUCT of mux21_8450 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25348
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25349
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25350
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8450
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8450 port map( A => n1, Y => n_S);
   NAND1 : nd2_25350 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25349 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25348 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8449 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8449;

architecture SYN_ARCHSTRUCT of mux21_8449 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25345
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25346
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25347
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8449
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8449 port map( A => n1, Y => n_S);
   NAND1 : nd2_25347 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25346 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25345 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8448 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8448;

architecture SYN_ARCHSTRUCT of mux21_8448 is

   component nd2_25342
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25343
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25344
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8448
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8448 port map( A => S, Y => n_S);
   NAND1 : nd2_25344 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25343 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25342 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8447 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8447;

architecture SYN_ARCHSTRUCT of mux21_8447 is

   component nd2_25339
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25340
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25341
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8447
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8447 port map( A => S, Y => n_S);
   NAND1 : nd2_25341 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25340 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25339 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8446 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8446;

architecture SYN_ARCHSTRUCT of mux21_8446 is

   component nd2_25336
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25337
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25338
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8446
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8446 port map( A => S, Y => n_S);
   NAND1 : nd2_25338 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25337 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25336 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8445 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8445;

architecture SYN_ARCHSTRUCT of mux21_8445 is

   component nd2_25333
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25334
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25335
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8445
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8445 port map( A => S, Y => n_S);
   NAND1 : nd2_25335 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25334 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25333 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8444 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8444;

architecture SYN_ARCHSTRUCT of mux21_8444 is

   component nd2_25330
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25331
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25332
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8444
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8444 port map( A => S, Y => n_S);
   NAND1 : nd2_25332 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25331 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25330 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8443 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8443;

architecture SYN_ARCHSTRUCT of mux21_8443 is

   component nd2_25327
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25328
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25329
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8443
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8443 port map( A => S, Y => n_S);
   NAND1 : nd2_25329 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25328 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25327 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8442 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8442;

architecture SYN_ARCHSTRUCT of mux21_8442 is

   component nd2_25324
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25325
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25326
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8442
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8442 port map( A => S, Y => n_S);
   NAND1 : nd2_25326 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25325 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25324 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8441 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8441;

architecture SYN_ARCHSTRUCT of mux21_8441 is

   component nd2_25321
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25322
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25323
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8441
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8441 port map( A => S, Y => n_S);
   NAND1 : nd2_25323 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25322 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25321 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8440 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8440;

architecture SYN_ARCHSTRUCT of mux21_8440 is

   component nd2_25318
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25319
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25320
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8440
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8440 port map( A => S, Y => n_S);
   NAND1 : nd2_25320 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25319 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25318 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8439 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8439;

architecture SYN_ARCHSTRUCT of mux21_8439 is

   component nd2_25315
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25316
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25317
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8439
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8439 port map( A => S, Y => n_S);
   NAND1 : nd2_25317 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25316 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25315 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8438 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8438;

architecture SYN_ARCHSTRUCT of mux21_8438 is

   component nd2_25312
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25313
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25314
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8438
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8438 port map( A => S, Y => n_S);
   NAND1 : nd2_25314 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25313 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25312 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8437 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8437;

architecture SYN_ARCHSTRUCT of mux21_8437 is

   component nd2_25309
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25310
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25311
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8437
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8437 port map( A => S, Y => n_S);
   NAND1 : nd2_25311 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25310 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25309 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8436 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8436;

architecture SYN_ARCHSTRUCT of mux21_8436 is

   component nd2_25306
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25307
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25308
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8436
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8436 port map( A => S, Y => n_S);
   NAND1 : nd2_25308 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25307 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25306 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8435 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8435;

architecture SYN_ARCHSTRUCT of mux21_8435 is

   component nd2_25303
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25304
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25305
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8435
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8435 port map( A => S, Y => n_S);
   NAND1 : nd2_25305 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25304 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25303 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8434 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8434;

architecture SYN_ARCHSTRUCT of mux21_8434 is

   component nd2_25300
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25301
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25302
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8434
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8434 port map( A => S, Y => n_S);
   NAND1 : nd2_25302 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25301 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25300 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8433 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8433;

architecture SYN_ARCHSTRUCT of mux21_8433 is

   component nd2_25297
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25298
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25299
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8433
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8433 port map( A => S, Y => n_S);
   NAND1 : nd2_25299 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25298 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25297 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8432 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8432;

architecture SYN_ARCHSTRUCT of mux21_8432 is

   component nd2_25294
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25295
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25296
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8432
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8432 port map( A => S, Y => n_S);
   NAND1 : nd2_25296 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25295 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25294 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8431 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8431;

architecture SYN_ARCHSTRUCT of mux21_8431 is

   component nd2_25291
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25292
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25293
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8431
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8431 port map( A => S, Y => n_S);
   NAND1 : nd2_25293 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25292 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25291 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8430 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8430;

architecture SYN_ARCHSTRUCT of mux21_8430 is

   component nd2_25288
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25289
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25290
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8430
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8430 port map( A => S, Y => n_S);
   NAND1 : nd2_25290 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25289 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25288 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8429 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8429;

architecture SYN_ARCHSTRUCT of mux21_8429 is

   component nd2_25285
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25286
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25287
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8429
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8429 port map( A => S, Y => n_S);
   NAND1 : nd2_25287 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25286 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25285 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8428 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8428;

architecture SYN_ARCHSTRUCT of mux21_8428 is

   component nd2_25282
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25283
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25284
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8428
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8428 port map( A => S, Y => n_S);
   NAND1 : nd2_25284 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25283 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25282 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8427 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8427;

architecture SYN_ARCHSTRUCT of mux21_8427 is

   component nd2_25279
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25280
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25281
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8427
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8427 port map( A => S, Y => n_S);
   NAND1 : nd2_25281 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25280 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25279 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8426 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8426;

architecture SYN_ARCHSTRUCT of mux21_8426 is

   component nd2_25276
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25277
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25278
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8426
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8426 port map( A => S, Y => n_S);
   NAND1 : nd2_25278 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25277 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25276 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8425 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8425;

architecture SYN_ARCHSTRUCT of mux21_8425 is

   component nd2_25273
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25274
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25275
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8425
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8425 port map( A => S, Y => n_S);
   NAND1 : nd2_25275 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25274 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25273 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8424 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8424;

architecture SYN_ARCHSTRUCT of mux21_8424 is

   component nd2_25270
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25271
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25272
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8424
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8424 port map( A => S, Y => n_S);
   NAND1 : nd2_25272 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25271 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25270 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8423 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8423;

architecture SYN_ARCHSTRUCT of mux21_8423 is

   component nd2_25267
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25268
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25269
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8423
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8423 port map( A => S, Y => n_S);
   NAND1 : nd2_25269 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25268 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25267 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8422 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8422;

architecture SYN_ARCHSTRUCT of mux21_8422 is

   component nd2_25264
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25265
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25266
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8422
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8422 port map( A => S, Y => n_S);
   NAND1 : nd2_25266 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25265 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25264 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8421 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8421;

architecture SYN_ARCHSTRUCT of mux21_8421 is

   component nd2_25261
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25262
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25263
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8421
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8421 port map( A => S, Y => n_S);
   NAND1 : nd2_25263 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25262 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25261 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8420 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8420;

architecture SYN_ARCHSTRUCT of mux21_8420 is

   component nd2_25258
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25259
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25260
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8420
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8420 port map( A => S, Y => n_S);
   NAND1 : nd2_25260 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25259 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25258 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8419 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8419;

architecture SYN_ARCHSTRUCT of mux21_8419 is

   component nd2_25255
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25256
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25257
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8419
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8419 port map( A => S, Y => n_S);
   NAND1 : nd2_25257 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25256 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25255 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8418 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8418;

architecture SYN_ARCHSTRUCT of mux21_8418 is

   component nd2_25252
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25253
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25254
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8418
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8418 port map( A => S, Y => n_S);
   NAND1 : nd2_25254 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25253 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25252 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8417 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8417;

architecture SYN_ARCHSTRUCT of mux21_8417 is

   component nd2_25249
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25250
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25251
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8417
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8417 port map( A => S, Y => n_S);
   NAND1 : nd2_25251 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25250 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25249 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8416 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8416;

architecture SYN_ARCHSTRUCT of mux21_8416 is

   component nd2_25246
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25247
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25248
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8416
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8416 port map( A => S, Y => n_S);
   NAND1 : nd2_25248 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25247 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25246 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8415 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8415;

architecture SYN_ARCHSTRUCT of mux21_8415 is

   component nd2_25243
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25244
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25245
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8415
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8415 port map( A => S, Y => n_S);
   NAND1 : nd2_25245 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25244 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25243 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8414 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8414;

architecture SYN_ARCHSTRUCT of mux21_8414 is

   component nd2_25240
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25241
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25242
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8414
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8414 port map( A => S, Y => n_S);
   NAND1 : nd2_25242 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25241 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25240 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8413 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8413;

architecture SYN_ARCHSTRUCT of mux21_8413 is

   component nd2_25237
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25238
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25239
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8413
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8413 port map( A => S, Y => n_S);
   NAND1 : nd2_25239 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25238 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25237 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8412 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8412;

architecture SYN_ARCHSTRUCT of mux21_8412 is

   component nd2_25234
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25235
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25236
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8412
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8412 port map( A => S, Y => n_S);
   NAND1 : nd2_25236 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25235 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25234 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8411 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8411;

architecture SYN_ARCHSTRUCT of mux21_8411 is

   component nd2_25231
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25232
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25233
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8411
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8411 port map( A => S, Y => n_S);
   NAND1 : nd2_25233 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25232 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25231 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8410 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8410;

architecture SYN_ARCHSTRUCT of mux21_8410 is

   component nd2_25228
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25229
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25230
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8410
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8410 port map( A => S, Y => n_S);
   NAND1 : nd2_25230 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25229 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25228 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8409 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8409;

architecture SYN_ARCHSTRUCT of mux21_8409 is

   component nd2_25225
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25226
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25227
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8409
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8409 port map( A => S, Y => n_S);
   NAND1 : nd2_25227 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25226 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25225 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8408 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8408;

architecture SYN_ARCHSTRUCT of mux21_8408 is

   component nd2_25222
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25223
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25224
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8408
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8408 port map( A => S, Y => n_S);
   NAND1 : nd2_25224 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25223 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25222 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8407 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8407;

architecture SYN_ARCHSTRUCT of mux21_8407 is

   component nd2_25219
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25220
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25221
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8407
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8407 port map( A => S, Y => n_S);
   NAND1 : nd2_25221 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25220 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25219 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8406 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8406;

architecture SYN_ARCHSTRUCT of mux21_8406 is

   component nd2_25216
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25217
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25218
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8406
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8406 port map( A => S, Y => n_S);
   NAND1 : nd2_25218 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25217 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25216 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8405 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8405;

architecture SYN_ARCHSTRUCT of mux21_8405 is

   component nd2_25213
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25214
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25215
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8405
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8405 port map( A => S, Y => n_S);
   NAND1 : nd2_25215 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25214 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25213 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8404 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8404;

architecture SYN_ARCHSTRUCT of mux21_8404 is

   component nd2_25210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25211
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25212
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8404
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8404 port map( A => S, Y => n_S);
   NAND1 : nd2_25212 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25211 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25210 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8403 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8403;

architecture SYN_ARCHSTRUCT of mux21_8403 is

   component nd2_25207
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25208
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25209
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8403
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8403 port map( A => S, Y => n_S);
   NAND1 : nd2_25209 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25208 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25207 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8402 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8402;

architecture SYN_ARCHSTRUCT of mux21_8402 is

   component nd2_25204
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25205
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25206
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8402
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8402 port map( A => S, Y => n_S);
   NAND1 : nd2_25206 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25205 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25204 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8401 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8401;

architecture SYN_ARCHSTRUCT of mux21_8401 is

   component nd2_25201
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25202
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25203
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8401
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8401 port map( A => S, Y => n_S);
   NAND1 : nd2_25203 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25202 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25201 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8400 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8400;

architecture SYN_ARCHSTRUCT of mux21_8400 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25198
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25199
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25200
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8400
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8400 port map( A => n1, Y => n_S);
   NAND1 : nd2_25200 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25199 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25198 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8399 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8399;

architecture SYN_ARCHSTRUCT of mux21_8399 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25195
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25196
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25197
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8399
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8399 port map( A => n1, Y => n_S);
   NAND1 : nd2_25197 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25196 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25195 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8398 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8398;

architecture SYN_ARCHSTRUCT of mux21_8398 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25192
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25193
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25194
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8398
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8398 port map( A => n1, Y => n_S);
   NAND1 : nd2_25194 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25193 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25192 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8397 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8397;

architecture SYN_ARCHSTRUCT of mux21_8397 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8397
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8397 port map( A => n1, Y => n_S);
   NAND1 : nd2_25191 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25190 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25189 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8396 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8396;

architecture SYN_ARCHSTRUCT of mux21_8396 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8396
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8396 port map( A => n1, Y => n_S);
   NAND1 : nd2_25188 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25187 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25186 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8395 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8395;

architecture SYN_ARCHSTRUCT of mux21_8395 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8395
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8395 port map( A => n1, Y => n_S);
   NAND1 : nd2_25185 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25184 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25183 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8394 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8394;

architecture SYN_ARCHSTRUCT of mux21_8394 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8394
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8394 port map( A => n1, Y => n_S);
   NAND1 : nd2_25182 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25181 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25180 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8393 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8393;

architecture SYN_ARCHSTRUCT of mux21_8393 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8393
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8393 port map( A => n1, Y => n_S);
   NAND1 : nd2_25179 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25178 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25177 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8392 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8392;

architecture SYN_ARCHSTRUCT of mux21_8392 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8392
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8392 port map( A => n1, Y => n_S);
   NAND1 : nd2_25176 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25175 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25174 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8391 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8391;

architecture SYN_ARCHSTRUCT of mux21_8391 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8391
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8391 port map( A => n1, Y => n_S);
   NAND1 : nd2_25173 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25172 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25171 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8390 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8390;

architecture SYN_ARCHSTRUCT of mux21_8390 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8390
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8390 port map( A => n1, Y => n_S);
   NAND1 : nd2_25170 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25169 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25168 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8389 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8389;

architecture SYN_ARCHSTRUCT of mux21_8389 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8389
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8389 port map( A => n1, Y => n_S);
   NAND1 : nd2_25167 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25166 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25165 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8388 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8388;

architecture SYN_ARCHSTRUCT of mux21_8388 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8388
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8388 port map( A => n1, Y => n_S);
   NAND1 : nd2_25164 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25163 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25162 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8387 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8387;

architecture SYN_ARCHSTRUCT of mux21_8387 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8387
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8387 port map( A => n1, Y => n_S);
   NAND1 : nd2_25161 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25160 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25159 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8386 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8386;

architecture SYN_ARCHSTRUCT of mux21_8386 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8386
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8386 port map( A => n1, Y => n_S);
   NAND1 : nd2_25158 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25157 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25156 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8385 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8385;

architecture SYN_ARCHSTRUCT of mux21_8385 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8385
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8385 port map( A => n1, Y => n_S);
   NAND1 : nd2_25155 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25154 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25153 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8384 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8384;

architecture SYN_ARCHSTRUCT of mux21_8384 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8384
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8384 port map( A => n1, Y => n_S);
   NAND1 : nd2_25152 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25151 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25150 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8383 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8383;

architecture SYN_ARCHSTRUCT of mux21_8383 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8383
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8383 port map( A => n1, Y => n_S);
   NAND1 : nd2_25149 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25148 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25147 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8382 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8382;

architecture SYN_ARCHSTRUCT of mux21_8382 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8382
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8382 port map( A => n1, Y => n_S);
   NAND1 : nd2_25146 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25145 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25144 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8381 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8381;

architecture SYN_ARCHSTRUCT of mux21_8381 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8381
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8381 port map( A => n1, Y => n_S);
   NAND1 : nd2_25143 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25142 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25141 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8380 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8380;

architecture SYN_ARCHSTRUCT of mux21_8380 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8380
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8380 port map( A => n1, Y => n_S);
   NAND1 : nd2_25140 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25139 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25138 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8379 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8379;

architecture SYN_ARCHSTRUCT of mux21_8379 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8379
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8379 port map( A => n1, Y => n_S);
   NAND1 : nd2_25137 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25136 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25135 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8378 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8378;

architecture SYN_ARCHSTRUCT of mux21_8378 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8378
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8378 port map( A => n1, Y => n_S);
   NAND1 : nd2_25134 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25133 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25132 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8377 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8377;

architecture SYN_ARCHSTRUCT of mux21_8377 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8377
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8377 port map( A => n1, Y => n_S);
   NAND1 : nd2_25131 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25130 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25129 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8376 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8376;

architecture SYN_ARCHSTRUCT of mux21_8376 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8376
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8376 port map( A => n1, Y => n_S);
   NAND1 : nd2_25128 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25127 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25126 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8375 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8375;

architecture SYN_ARCHSTRUCT of mux21_8375 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8375
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8375 port map( A => n1, Y => n_S);
   NAND1 : nd2_25125 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25124 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25123 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8374 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8374;

architecture SYN_ARCHSTRUCT of mux21_8374 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8374
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8374 port map( A => n1, Y => n_S);
   NAND1 : nd2_25122 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25121 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25120 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8373 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8373;

architecture SYN_ARCHSTRUCT of mux21_8373 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8373
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8373 port map( A => n1, Y => n_S);
   NAND1 : nd2_25119 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25118 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25117 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8372 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8372;

architecture SYN_ARCHSTRUCT of mux21_8372 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8372
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8372 port map( A => n1, Y => n_S);
   NAND1 : nd2_25116 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25115 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25114 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8371 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8371;

architecture SYN_ARCHSTRUCT of mux21_8371 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8371
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8371 port map( A => n1, Y => n_S);
   NAND1 : nd2_25113 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25112 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25111 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8370 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8370;

architecture SYN_ARCHSTRUCT of mux21_8370 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8370
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8370 port map( A => n1, Y => n_S);
   NAND1 : nd2_25110 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25109 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25108 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8369 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8369;

architecture SYN_ARCHSTRUCT of mux21_8369 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8369
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8369 port map( A => n1, Y => n_S);
   NAND1 : nd2_25107 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25106 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25105 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8368 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8368;

architecture SYN_ARCHSTRUCT of mux21_8368 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8368
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8368 port map( A => n1, Y => n_S);
   NAND1 : nd2_25104 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25103 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25102 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8367 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8367;

architecture SYN_ARCHSTRUCT of mux21_8367 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25099
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8367
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8367 port map( A => n1, Y => n_S);
   NAND1 : nd2_25101 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25100 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25099 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8366 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8366;

architecture SYN_ARCHSTRUCT of mux21_8366 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25096
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25097
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25098
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8366
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8366 port map( A => n1, Y => n_S);
   NAND1 : nd2_25098 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25097 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25096 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8365 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8365;

architecture SYN_ARCHSTRUCT of mux21_8365 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25093
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25094
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25095
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8365
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8365 port map( A => n1, Y => n_S);
   NAND1 : nd2_25095 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25094 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25093 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8364 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8364;

architecture SYN_ARCHSTRUCT of mux21_8364 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25090
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25091
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25092
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8364
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8364 port map( A => n1, Y => n_S);
   NAND1 : nd2_25092 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25091 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25090 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8363 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8363;

architecture SYN_ARCHSTRUCT of mux21_8363 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25087
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25088
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25089
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8363
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8363 port map( A => n1, Y => n_S);
   NAND1 : nd2_25089 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25088 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25087 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8362 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8362;

architecture SYN_ARCHSTRUCT of mux21_8362 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25084
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25085
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25086
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8362
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8362 port map( A => n1, Y => n_S);
   NAND1 : nd2_25086 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25085 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25084 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8361 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8361;

architecture SYN_ARCHSTRUCT of mux21_8361 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25081
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25082
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25083
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8361
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8361 port map( A => n1, Y => n_S);
   NAND1 : nd2_25083 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25082 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25081 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8360 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8360;

architecture SYN_ARCHSTRUCT of mux21_8360 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25078
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25079
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25080
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8360
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8360 port map( A => n1, Y => n_S);
   NAND1 : nd2_25080 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25079 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25078 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8359 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8359;

architecture SYN_ARCHSTRUCT of mux21_8359 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25075
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25076
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25077
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8359
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8359 port map( A => n1, Y => n_S);
   NAND1 : nd2_25077 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25076 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25075 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8358 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8358;

architecture SYN_ARCHSTRUCT of mux21_8358 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25072
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25073
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25074
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8358
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8358 port map( A => n1, Y => n_S);
   NAND1 : nd2_25074 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25073 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25072 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8357 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8357;

architecture SYN_ARCHSTRUCT of mux21_8357 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25069
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25070
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25071
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8357
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8357 port map( A => n1, Y => n_S);
   NAND1 : nd2_25071 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25070 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25069 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8356 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8356;

architecture SYN_ARCHSTRUCT of mux21_8356 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25066
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25067
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25068
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8356
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8356 port map( A => n1, Y => n_S);
   NAND1 : nd2_25068 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25067 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25066 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8355 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8355;

architecture SYN_ARCHSTRUCT of mux21_8355 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25063
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25064
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25065
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8355
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8355 port map( A => n1, Y => n_S);
   NAND1 : nd2_25065 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25064 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25063 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8354 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8354;

architecture SYN_ARCHSTRUCT of mux21_8354 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25060
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25061
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25062
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8354
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8354 port map( A => n1, Y => n_S);
   NAND1 : nd2_25062 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25061 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25060 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8353 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8353;

architecture SYN_ARCHSTRUCT of mux21_8353 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25057
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25058
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25059
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8353
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8353 port map( A => n1, Y => n_S);
   NAND1 : nd2_25059 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25058 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25057 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8352 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8352;

architecture SYN_ARCHSTRUCT of mux21_8352 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25054
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25055
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25056
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8352
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8352 port map( A => n1, Y => n_S);
   NAND1 : nd2_25056 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25055 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25054 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8351 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8351;

architecture SYN_ARCHSTRUCT of mux21_8351 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25051
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25052
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25053
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8351
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8351 port map( A => n1, Y => n_S);
   NAND1 : nd2_25053 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25052 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25051 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8350 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8350;

architecture SYN_ARCHSTRUCT of mux21_8350 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25048
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25049
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25050
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8350
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8350 port map( A => n1, Y => n_S);
   NAND1 : nd2_25050 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25049 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25048 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8349 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8349;

architecture SYN_ARCHSTRUCT of mux21_8349 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25045
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25046
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25047
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8349
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8349 port map( A => n1, Y => n_S);
   NAND1 : nd2_25047 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25046 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25045 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8348 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8348;

architecture SYN_ARCHSTRUCT of mux21_8348 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25042
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25043
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25044
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8348
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8348 port map( A => n1, Y => n_S);
   NAND1 : nd2_25044 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25043 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25042 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8347 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8347;

architecture SYN_ARCHSTRUCT of mux21_8347 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25039
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25040
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25041
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8347
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8347 port map( A => n1, Y => n_S);
   NAND1 : nd2_25041 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25040 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25039 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8346 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8346;

architecture SYN_ARCHSTRUCT of mux21_8346 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25036
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25037
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25038
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8346
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8346 port map( A => n1, Y => n_S);
   NAND1 : nd2_25038 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25037 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25036 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8345 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8345;

architecture SYN_ARCHSTRUCT of mux21_8345 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25033
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25034
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25035
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8345
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8345 port map( A => n1, Y => n_S);
   NAND1 : nd2_25035 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25034 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25033 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8344 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8344;

architecture SYN_ARCHSTRUCT of mux21_8344 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25030
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25031
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25032
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8344
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8344 port map( A => n1, Y => n_S);
   NAND1 : nd2_25032 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25031 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25030 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8343 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8343;

architecture SYN_ARCHSTRUCT of mux21_8343 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25027
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25028
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25029
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8343
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8343 port map( A => n1, Y => n_S);
   NAND1 : nd2_25029 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25028 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25027 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8342 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8342;

architecture SYN_ARCHSTRUCT of mux21_8342 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25024
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25025
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25026
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8342
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8342 port map( A => n1, Y => n_S);
   NAND1 : nd2_25026 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25025 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25024 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8341 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8341;

architecture SYN_ARCHSTRUCT of mux21_8341 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25021
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25022
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25023
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8341
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8341 port map( A => n1, Y => n_S);
   NAND1 : nd2_25023 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25022 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25021 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8340 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8340;

architecture SYN_ARCHSTRUCT of mux21_8340 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25018
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25019
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25020
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8340
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8340 port map( A => n1, Y => n_S);
   NAND1 : nd2_25020 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25019 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25018 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8339 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8339;

architecture SYN_ARCHSTRUCT of mux21_8339 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25015
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25016
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25017
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8339
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8339 port map( A => n1, Y => n_S);
   NAND1 : nd2_25017 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25016 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25015 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8338 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8338;

architecture SYN_ARCHSTRUCT of mux21_8338 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25012
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25013
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25014
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8338
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8338 port map( A => n1, Y => n_S);
   NAND1 : nd2_25014 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25013 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25012 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8337 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8337;

architecture SYN_ARCHSTRUCT of mux21_8337 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25009
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25010
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25011
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8337
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8337 port map( A => n1, Y => n_S);
   NAND1 : nd2_25011 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25010 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25009 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8336 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8336;

architecture SYN_ARCHSTRUCT of mux21_8336 is

   component nd2_25006
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25007
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25008
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8336
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8336 port map( A => S, Y => n_S);
   NAND1 : nd2_25008 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25007 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25006 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8335 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8335;

architecture SYN_ARCHSTRUCT of mux21_8335 is

   component nd2_25003
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25004
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25005
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8335
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8335 port map( A => S, Y => n_S);
   NAND1 : nd2_25005 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25004 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25003 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8334 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8334;

architecture SYN_ARCHSTRUCT of mux21_8334 is

   component nd2_25000
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25001
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25002
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8334
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8334 port map( A => S, Y => n_S);
   NAND1 : nd2_25002 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_25001 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25000 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8333 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8333;

architecture SYN_ARCHSTRUCT of mux21_8333 is

   component nd2_24997
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24998
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24999
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8333
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8333 port map( A => S, Y => n_S);
   NAND1 : nd2_24999 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24998 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24997 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8332 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8332;

architecture SYN_ARCHSTRUCT of mux21_8332 is

   component nd2_24994
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24995
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24996
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8332
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8332 port map( A => S, Y => n_S);
   NAND1 : nd2_24996 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24995 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24994 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8331 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8331;

architecture SYN_ARCHSTRUCT of mux21_8331 is

   component nd2_24991
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24992
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24993
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8331
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8331 port map( A => S, Y => n_S);
   NAND1 : nd2_24993 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24992 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24991 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8330 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8330;

architecture SYN_ARCHSTRUCT of mux21_8330 is

   component nd2_24988
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24989
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24990
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8330
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8330 port map( A => S, Y => n_S);
   NAND1 : nd2_24990 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24989 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24988 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8329 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8329;

architecture SYN_ARCHSTRUCT of mux21_8329 is

   component nd2_24985
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24986
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24987
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8329
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8329 port map( A => S, Y => n_S);
   NAND1 : nd2_24987 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24986 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24985 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8328 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8328;

architecture SYN_ARCHSTRUCT of mux21_8328 is

   component nd2_24982
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24983
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24984
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8328
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8328 port map( A => S, Y => n_S);
   NAND1 : nd2_24984 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24983 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24982 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8327 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8327;

architecture SYN_ARCHSTRUCT of mux21_8327 is

   component nd2_24979
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24980
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24981
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8327
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8327 port map( A => S, Y => n_S);
   NAND1 : nd2_24981 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24980 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24979 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8326 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8326;

architecture SYN_ARCHSTRUCT of mux21_8326 is

   component nd2_24976
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24977
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24978
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8326
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8326 port map( A => S, Y => n_S);
   NAND1 : nd2_24978 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24977 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24976 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8325 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8325;

architecture SYN_ARCHSTRUCT of mux21_8325 is

   component nd2_24973
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24974
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24975
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8325
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8325 port map( A => S, Y => n_S);
   NAND1 : nd2_24975 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24974 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24973 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8324 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8324;

architecture SYN_ARCHSTRUCT of mux21_8324 is

   component nd2_24970
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24971
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24972
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8324
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8324 port map( A => S, Y => n_S);
   NAND1 : nd2_24972 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24971 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24970 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8323 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8323;

architecture SYN_ARCHSTRUCT of mux21_8323 is

   component nd2_24967
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24968
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24969
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8323
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8323 port map( A => S, Y => n_S);
   NAND1 : nd2_24969 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24968 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24967 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8322 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8322;

architecture SYN_ARCHSTRUCT of mux21_8322 is

   component nd2_24964
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24965
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24966
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8322
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8322 port map( A => S, Y => n_S);
   NAND1 : nd2_24966 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24965 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24964 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8321 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8321;

architecture SYN_ARCHSTRUCT of mux21_8321 is

   component nd2_24961
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24962
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24963
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8321
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8321 port map( A => S, Y => n_S);
   NAND1 : nd2_24963 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24962 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24961 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8320 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8320;

architecture SYN_ARCHSTRUCT of mux21_8320 is

   component nd2_24958
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24959
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24960
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8320
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8320 port map( A => S, Y => n_S);
   NAND1 : nd2_24960 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24959 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24958 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8319 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8319;

architecture SYN_ARCHSTRUCT of mux21_8319 is

   component nd2_24955
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24956
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24957
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8319
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8319 port map( A => S, Y => n_S);
   NAND1 : nd2_24957 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24956 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24955 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8318 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8318;

architecture SYN_ARCHSTRUCT of mux21_8318 is

   component nd2_24952
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24953
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24954
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8318
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8318 port map( A => S, Y => n_S);
   NAND1 : nd2_24954 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24953 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24952 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8317 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8317;

architecture SYN_ARCHSTRUCT of mux21_8317 is

   component nd2_24949
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24950
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24951
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8317
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8317 port map( A => S, Y => n_S);
   NAND1 : nd2_24951 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24950 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24949 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8316 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8316;

architecture SYN_ARCHSTRUCT of mux21_8316 is

   component nd2_24946
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24947
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24948
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8316
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8316 port map( A => S, Y => n_S);
   NAND1 : nd2_24948 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24947 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24946 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8315 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8315;

architecture SYN_ARCHSTRUCT of mux21_8315 is

   component nd2_24943
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24944
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24945
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8315
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8315 port map( A => S, Y => n_S);
   NAND1 : nd2_24945 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24944 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24943 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8314 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8314;

architecture SYN_ARCHSTRUCT of mux21_8314 is

   component nd2_24940
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24941
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24942
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8314
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8314 port map( A => S, Y => n_S);
   NAND1 : nd2_24942 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24941 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24940 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8313 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8313;

architecture SYN_ARCHSTRUCT of mux21_8313 is

   component nd2_24937
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24938
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24939
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8313
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8313 port map( A => S, Y => n_S);
   NAND1 : nd2_24939 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24938 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24937 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8312 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8312;

architecture SYN_ARCHSTRUCT of mux21_8312 is

   component nd2_24934
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24935
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24936
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8312
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8312 port map( A => S, Y => n_S);
   NAND1 : nd2_24936 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24935 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24934 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8311 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8311;

architecture SYN_ARCHSTRUCT of mux21_8311 is

   component nd2_24931
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24932
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24933
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8311
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8311 port map( A => S, Y => n_S);
   NAND1 : nd2_24933 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24932 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24931 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8310 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8310;

architecture SYN_ARCHSTRUCT of mux21_8310 is

   component nd2_24928
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24929
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24930
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8310
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8310 port map( A => S, Y => n_S);
   NAND1 : nd2_24930 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24929 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24928 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8309 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8309;

architecture SYN_ARCHSTRUCT of mux21_8309 is

   component nd2_24925
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24926
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24927
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8309
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8309 port map( A => S, Y => n_S);
   NAND1 : nd2_24927 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24926 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24925 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8308 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8308;

architecture SYN_ARCHSTRUCT of mux21_8308 is

   component nd2_24922
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24923
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24924
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8308
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8308 port map( A => S, Y => n_S);
   NAND1 : nd2_24924 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24923 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24922 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8307 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8307;

architecture SYN_ARCHSTRUCT of mux21_8307 is

   component nd2_24919
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24920
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24921
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8307
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8307 port map( A => S, Y => n_S);
   NAND1 : nd2_24921 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24920 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24919 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8306 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8306;

architecture SYN_ARCHSTRUCT of mux21_8306 is

   component nd2_24916
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24917
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24918
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8306
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8306 port map( A => S, Y => n_S);
   NAND1 : nd2_24918 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24917 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24916 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8305 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8305;

architecture SYN_ARCHSTRUCT of mux21_8305 is

   component nd2_24913
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24914
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24915
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8305
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8305 port map( A => S, Y => n_S);
   NAND1 : nd2_24915 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24914 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24913 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8304 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8304;

architecture SYN_ARCHSTRUCT of mux21_8304 is

   component nd2_24910
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24911
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24912
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8304
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8304 port map( A => S, Y => n_S);
   NAND1 : nd2_24912 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24911 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24910 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8303 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8303;

architecture SYN_ARCHSTRUCT of mux21_8303 is

   component nd2_24907
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24908
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24909
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8303
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8303 port map( A => S, Y => n_S);
   NAND1 : nd2_24909 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24908 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24907 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8302 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8302;

architecture SYN_ARCHSTRUCT of mux21_8302 is

   component nd2_24904
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24905
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24906
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8302
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8302 port map( A => S, Y => n_S);
   NAND1 : nd2_24906 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24905 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24904 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8301 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8301;

architecture SYN_ARCHSTRUCT of mux21_8301 is

   component nd2_24901
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24902
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24903
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8301
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8301 port map( A => S, Y => n_S);
   NAND1 : nd2_24903 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24902 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24901 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8300 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8300;

architecture SYN_ARCHSTRUCT of mux21_8300 is

   component nd2_24898
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24899
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24900
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8300
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8300 port map( A => S, Y => n_S);
   NAND1 : nd2_24900 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24899 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24898 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8299 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8299;

architecture SYN_ARCHSTRUCT of mux21_8299 is

   component nd2_24895
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24896
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24897
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8299
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8299 port map( A => S, Y => n_S);
   NAND1 : nd2_24897 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24896 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24895 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8298 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8298;

architecture SYN_ARCHSTRUCT of mux21_8298 is

   component nd2_24892
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24893
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24894
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8298
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8298 port map( A => S, Y => n_S);
   NAND1 : nd2_24894 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24893 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24892 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8297 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8297;

architecture SYN_ARCHSTRUCT of mux21_8297 is

   component nd2_24889
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24890
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24891
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8297
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8297 port map( A => S, Y => n_S);
   NAND1 : nd2_24891 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24890 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24889 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8296 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8296;

architecture SYN_ARCHSTRUCT of mux21_8296 is

   component nd2_24886
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24887
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24888
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8296
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8296 port map( A => S, Y => n_S);
   NAND1 : nd2_24888 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24887 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24886 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8295 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8295;

architecture SYN_ARCHSTRUCT of mux21_8295 is

   component nd2_24883
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24884
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24885
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8295
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8295 port map( A => S, Y => n_S);
   NAND1 : nd2_24885 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24884 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24883 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8294 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8294;

architecture SYN_ARCHSTRUCT of mux21_8294 is

   component nd2_24880
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24881
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24882
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8294
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8294 port map( A => S, Y => n_S);
   NAND1 : nd2_24882 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24881 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24880 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8293 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8293;

architecture SYN_ARCHSTRUCT of mux21_8293 is

   component nd2_24877
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24878
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24879
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8293
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8293 port map( A => S, Y => n_S);
   NAND1 : nd2_24879 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24878 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24877 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8292 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8292;

architecture SYN_ARCHSTRUCT of mux21_8292 is

   component nd2_24874
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24875
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24876
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8292
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8292 port map( A => S, Y => n_S);
   NAND1 : nd2_24876 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24875 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24874 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8291 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8291;

architecture SYN_ARCHSTRUCT of mux21_8291 is

   component nd2_24871
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24872
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24873
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8291
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8291 port map( A => S, Y => n_S);
   NAND1 : nd2_24873 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24872 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24871 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8290 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8290;

architecture SYN_ARCHSTRUCT of mux21_8290 is

   component nd2_24868
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24869
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24870
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8290
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8290 port map( A => S, Y => n_S);
   NAND1 : nd2_24870 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24869 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24868 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8289 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8289;

architecture SYN_ARCHSTRUCT of mux21_8289 is

   component nd2_24865
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24866
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24867
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8289
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8289 port map( A => S, Y => n_S);
   NAND1 : nd2_24867 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24866 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24865 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8288 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8288;

architecture SYN_ARCHSTRUCT of mux21_8288 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24862
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24863
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24864
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8288
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8288 port map( A => n1, Y => n_S);
   NAND1 : nd2_24864 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24863 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24862 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8287 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8287;

architecture SYN_ARCHSTRUCT of mux21_8287 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24859
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24860
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24861
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8287
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8287 port map( A => n1, Y => n_S);
   NAND1 : nd2_24861 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24860 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24859 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8286 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8286;

architecture SYN_ARCHSTRUCT of mux21_8286 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24856
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24857
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24858
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8286
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8286 port map( A => n1, Y => n_S);
   NAND1 : nd2_24858 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24857 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24856 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8285 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8285;

architecture SYN_ARCHSTRUCT of mux21_8285 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24853
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24854
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24855
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8285
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8285 port map( A => n1, Y => n_S);
   NAND1 : nd2_24855 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24854 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24853 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8284 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8284;

architecture SYN_ARCHSTRUCT of mux21_8284 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24850
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24851
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24852
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8284
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8284 port map( A => n1, Y => n_S);
   NAND1 : nd2_24852 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24851 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24850 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8283 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8283;

architecture SYN_ARCHSTRUCT of mux21_8283 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24847
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24848
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24849
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8283
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8283 port map( A => n1, Y => n_S);
   NAND1 : nd2_24849 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24848 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24847 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8282 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8282;

architecture SYN_ARCHSTRUCT of mux21_8282 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24844
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24845
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24846
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8282
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8282 port map( A => n1, Y => n_S);
   NAND1 : nd2_24846 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24845 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24844 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8281 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8281;

architecture SYN_ARCHSTRUCT of mux21_8281 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24841
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24842
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24843
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8281
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8281 port map( A => n1, Y => n_S);
   NAND1 : nd2_24843 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24842 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24841 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8280 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8280;

architecture SYN_ARCHSTRUCT of mux21_8280 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24838
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24839
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24840
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8280
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8280 port map( A => n1, Y => n_S);
   NAND1 : nd2_24840 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24839 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24838 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8279 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8279;

architecture SYN_ARCHSTRUCT of mux21_8279 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24835
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24836
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24837
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8279
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8279 port map( A => n1, Y => n_S);
   NAND1 : nd2_24837 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24836 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24835 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8278 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8278;

architecture SYN_ARCHSTRUCT of mux21_8278 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24832
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24833
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24834
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8278
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8278 port map( A => n1, Y => n_S);
   NAND1 : nd2_24834 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24833 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24832 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8277 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8277;

architecture SYN_ARCHSTRUCT of mux21_8277 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24829
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24830
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24831
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8277
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8277 port map( A => n1, Y => n_S);
   NAND1 : nd2_24831 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24830 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24829 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8276 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8276;

architecture SYN_ARCHSTRUCT of mux21_8276 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24826
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24827
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24828
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8276
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8276 port map( A => n1, Y => n_S);
   NAND1 : nd2_24828 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24827 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24826 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8275 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8275;

architecture SYN_ARCHSTRUCT of mux21_8275 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24823
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24824
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24825
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8275
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8275 port map( A => n1, Y => n_S);
   NAND1 : nd2_24825 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24824 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24823 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8274 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8274;

architecture SYN_ARCHSTRUCT of mux21_8274 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24820
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24821
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24822
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8274
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8274 port map( A => n1, Y => n_S);
   NAND1 : nd2_24822 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24821 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24820 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8273 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8273;

architecture SYN_ARCHSTRUCT of mux21_8273 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24817
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24818
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24819
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8273
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8273 port map( A => n1, Y => n_S);
   NAND1 : nd2_24819 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24818 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24817 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8272 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8272;

architecture SYN_ARCHSTRUCT of mux21_8272 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24814
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24815
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24816
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8272
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8272 port map( A => n1, Y => n_S);
   NAND1 : nd2_24816 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24815 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24814 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8271 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8271;

architecture SYN_ARCHSTRUCT of mux21_8271 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24811
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24812
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24813
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8271
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8271 port map( A => n1, Y => n_S);
   NAND1 : nd2_24813 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24812 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24811 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8270 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8270;

architecture SYN_ARCHSTRUCT of mux21_8270 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24808
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24809
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24810
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8270
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8270 port map( A => n1, Y => n_S);
   NAND1 : nd2_24810 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24809 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24808 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8269 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8269;

architecture SYN_ARCHSTRUCT of mux21_8269 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24805
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24806
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24807
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8269
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8269 port map( A => n1, Y => n_S);
   NAND1 : nd2_24807 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24806 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24805 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8268 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8268;

architecture SYN_ARCHSTRUCT of mux21_8268 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24802
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24803
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24804
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8268
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8268 port map( A => n1, Y => n_S);
   NAND1 : nd2_24804 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24803 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24802 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8267 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8267;

architecture SYN_ARCHSTRUCT of mux21_8267 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24799
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24800
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24801
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8267
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8267 port map( A => n1, Y => n_S);
   NAND1 : nd2_24801 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24800 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24799 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8266 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8266;

architecture SYN_ARCHSTRUCT of mux21_8266 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24796
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24797
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24798
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8266
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8266 port map( A => n1, Y => n_S);
   NAND1 : nd2_24798 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24797 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24796 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8265 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8265;

architecture SYN_ARCHSTRUCT of mux21_8265 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24793
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24794
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24795
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8265
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8265 port map( A => n1, Y => n_S);
   NAND1 : nd2_24795 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24794 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24793 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8264 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8264;

architecture SYN_ARCHSTRUCT of mux21_8264 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24790
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24791
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24792
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8264
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8264 port map( A => n1, Y => n_S);
   NAND1 : nd2_24792 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24791 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24790 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8263 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8263;

architecture SYN_ARCHSTRUCT of mux21_8263 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24787
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24788
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24789
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8263
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8263 port map( A => n1, Y => n_S);
   NAND1 : nd2_24789 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24788 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24787 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8262 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8262;

architecture SYN_ARCHSTRUCT of mux21_8262 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24784
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24785
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24786
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8262
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8262 port map( A => n1, Y => n_S);
   NAND1 : nd2_24786 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24785 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24784 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8261 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8261;

architecture SYN_ARCHSTRUCT of mux21_8261 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24781
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24782
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24783
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8261
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8261 port map( A => n1, Y => n_S);
   NAND1 : nd2_24783 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24782 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24781 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8260 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8260;

architecture SYN_ARCHSTRUCT of mux21_8260 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24778
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24779
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24780
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8260
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8260 port map( A => n1, Y => n_S);
   NAND1 : nd2_24780 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24779 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24778 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8259 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8259;

architecture SYN_ARCHSTRUCT of mux21_8259 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24775
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24776
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24777
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8259
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8259 port map( A => n1, Y => n_S);
   NAND1 : nd2_24777 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24776 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24775 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8258 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8258;

architecture SYN_ARCHSTRUCT of mux21_8258 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24772
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24773
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24774
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8258
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8258 port map( A => n1, Y => n_S);
   NAND1 : nd2_24774 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24773 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24772 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8257 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8257;

architecture SYN_ARCHSTRUCT of mux21_8257 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24769
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24770
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24771
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8257
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8257 port map( A => n1, Y => n_S);
   NAND1 : nd2_24771 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24770 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24769 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8256 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8256;

architecture SYN_ARCHSTRUCT of mux21_8256 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24766
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24767
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24768
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8256
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8256 port map( A => n1, Y => n_S);
   NAND1 : nd2_24768 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24767 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24766 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8255 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8255;

architecture SYN_ARCHSTRUCT of mux21_8255 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24763
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24764
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24765
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8255
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8255 port map( A => n1, Y => n_S);
   NAND1 : nd2_24765 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24764 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24763 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8254 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8254;

architecture SYN_ARCHSTRUCT of mux21_8254 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24760
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24761
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24762
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8254
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8254 port map( A => n1, Y => n_S);
   NAND1 : nd2_24762 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24761 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24760 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8253 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8253;

architecture SYN_ARCHSTRUCT of mux21_8253 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24757
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24758
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24759
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8253
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8253 port map( A => n1, Y => n_S);
   NAND1 : nd2_24759 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24758 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24757 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8252 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8252;

architecture SYN_ARCHSTRUCT of mux21_8252 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24754
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24755
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24756
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8252
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8252 port map( A => n1, Y => n_S);
   NAND1 : nd2_24756 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24755 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24754 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8251 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8251;

architecture SYN_ARCHSTRUCT of mux21_8251 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24751
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24752
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24753
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8251
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8251 port map( A => n1, Y => n_S);
   NAND1 : nd2_24753 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24752 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24751 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8250 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8250;

architecture SYN_ARCHSTRUCT of mux21_8250 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24748
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24749
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24750
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8250
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8250 port map( A => n1, Y => n_S);
   NAND1 : nd2_24750 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24749 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24748 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8249 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8249;

architecture SYN_ARCHSTRUCT of mux21_8249 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24745
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24746
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24747
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8249
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8249 port map( A => n1, Y => n_S);
   NAND1 : nd2_24747 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24746 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24745 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8248 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8248;

architecture SYN_ARCHSTRUCT of mux21_8248 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24742
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24743
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24744
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8248
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8248 port map( A => n1, Y => n_S);
   NAND1 : nd2_24744 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24743 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24742 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8247 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8247;

architecture SYN_ARCHSTRUCT of mux21_8247 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24739
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24740
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24741
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8247
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8247 port map( A => n1, Y => n_S);
   NAND1 : nd2_24741 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24740 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24739 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8246 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8246;

architecture SYN_ARCHSTRUCT of mux21_8246 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24736
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24737
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24738
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8246
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8246 port map( A => n1, Y => n_S);
   NAND1 : nd2_24738 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24737 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24736 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8245 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8245;

architecture SYN_ARCHSTRUCT of mux21_8245 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24733
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24734
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24735
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8245
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8245 port map( A => n1, Y => n_S);
   NAND1 : nd2_24735 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24734 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24733 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8244 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8244;

architecture SYN_ARCHSTRUCT of mux21_8244 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24730
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24731
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24732
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8244
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8244 port map( A => n1, Y => n_S);
   NAND1 : nd2_24732 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24731 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24730 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8243 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8243;

architecture SYN_ARCHSTRUCT of mux21_8243 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24727
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24728
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24729
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8243
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8243 port map( A => n1, Y => n_S);
   NAND1 : nd2_24729 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24728 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24727 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8242 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8242;

architecture SYN_ARCHSTRUCT of mux21_8242 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24724
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24725
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24726
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8242
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8242 port map( A => n1, Y => n_S);
   NAND1 : nd2_24726 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24725 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24724 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8241 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8241;

architecture SYN_ARCHSTRUCT of mux21_8241 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24721
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24722
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24723
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8241
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8241 port map( A => n1, Y => n_S);
   NAND1 : nd2_24723 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24722 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24721 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8240 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8240;

architecture SYN_ARCHSTRUCT of mux21_8240 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24718
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24719
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24720
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8240
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8240 port map( A => n1, Y => n_S);
   NAND1 : nd2_24720 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24719 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24718 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8239 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8239;

architecture SYN_ARCHSTRUCT of mux21_8239 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24715
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24716
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24717
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8239
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8239 port map( A => n1, Y => n_S);
   NAND1 : nd2_24717 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24716 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24715 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8238 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8238;

architecture SYN_ARCHSTRUCT of mux21_8238 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24712
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24713
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24714
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8238
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8238 port map( A => n1, Y => n_S);
   NAND1 : nd2_24714 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24713 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24712 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8237 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8237;

architecture SYN_ARCHSTRUCT of mux21_8237 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24709
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24710
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24711
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8237
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8237 port map( A => n1, Y => n_S);
   NAND1 : nd2_24711 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24710 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24709 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8236 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8236;

architecture SYN_ARCHSTRUCT of mux21_8236 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24706
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24707
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24708
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8236
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8236 port map( A => n1, Y => n_S);
   NAND1 : nd2_24708 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24707 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24706 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8235 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8235;

architecture SYN_ARCHSTRUCT of mux21_8235 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24703
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24704
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24705
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8235
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8235 port map( A => n1, Y => n_S);
   NAND1 : nd2_24705 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24704 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24703 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8234 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8234;

architecture SYN_ARCHSTRUCT of mux21_8234 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24700
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24701
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24702
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8234
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8234 port map( A => n1, Y => n_S);
   NAND1 : nd2_24702 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24701 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24700 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8233 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8233;

architecture SYN_ARCHSTRUCT of mux21_8233 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24697
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24698
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24699
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8233
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8233 port map( A => n1, Y => n_S);
   NAND1 : nd2_24699 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24698 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24697 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8232 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8232;

architecture SYN_ARCHSTRUCT of mux21_8232 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24694
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24695
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24696
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8232
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8232 port map( A => n1, Y => n_S);
   NAND1 : nd2_24696 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24695 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24694 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8231 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8231;

architecture SYN_ARCHSTRUCT of mux21_8231 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24691
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24692
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24693
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8231
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8231 port map( A => n1, Y => n_S);
   NAND1 : nd2_24693 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24692 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24691 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8230 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8230;

architecture SYN_ARCHSTRUCT of mux21_8230 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24688
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24689
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24690
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8230
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8230 port map( A => n1, Y => n_S);
   NAND1 : nd2_24690 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24689 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24688 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8229 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8229;

architecture SYN_ARCHSTRUCT of mux21_8229 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24685
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24686
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24687
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8229
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8229 port map( A => n1, Y => n_S);
   NAND1 : nd2_24687 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24686 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24685 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8228 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8228;

architecture SYN_ARCHSTRUCT of mux21_8228 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24682
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24683
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24684
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8228
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8228 port map( A => n1, Y => n_S);
   NAND1 : nd2_24684 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24683 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24682 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8227 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8227;

architecture SYN_ARCHSTRUCT of mux21_8227 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24679
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24680
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24681
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8227
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8227 port map( A => n1, Y => n_S);
   NAND1 : nd2_24681 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24680 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24679 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8226 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8226;

architecture SYN_ARCHSTRUCT of mux21_8226 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24676
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24677
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24678
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8226
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8226 port map( A => n1, Y => n_S);
   NAND1 : nd2_24678 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24677 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24676 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8225 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8225;

architecture SYN_ARCHSTRUCT of mux21_8225 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_24673
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24674
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24675
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8225
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8225 port map( A => n1, Y => n_S);
   NAND1 : nd2_24675 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_24674 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24673 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8224 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8224;

architecture SYN_ARCHSTRUCT of mux21_8224 is

   component nd2_24670
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24671
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24672
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8224
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8224 port map( A => S, Y => n_S);
   NAND1 : nd2_24672 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24671 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24670 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8223 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8223;

architecture SYN_ARCHSTRUCT of mux21_8223 is

   component nd2_24667
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24668
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24669
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8223
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8223 port map( A => S, Y => n_S);
   NAND1 : nd2_24669 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24668 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24667 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8222 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8222;

architecture SYN_ARCHSTRUCT of mux21_8222 is

   component nd2_24664
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24665
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24666
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8222
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8222 port map( A => S, Y => n_S);
   NAND1 : nd2_24666 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24665 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24664 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8221 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8221;

architecture SYN_ARCHSTRUCT of mux21_8221 is

   component nd2_24661
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24662
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24663
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8221
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8221 port map( A => S, Y => n_S);
   NAND1 : nd2_24663 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24662 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24661 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8220 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8220;

architecture SYN_ARCHSTRUCT of mux21_8220 is

   component nd2_24658
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24659
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24660
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8220
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8220 port map( A => S, Y => n_S);
   NAND1 : nd2_24660 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24659 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24658 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8219 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8219;

architecture SYN_ARCHSTRUCT of mux21_8219 is

   component nd2_24655
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24656
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24657
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8219
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8219 port map( A => S, Y => n_S);
   NAND1 : nd2_24657 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24656 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24655 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8218 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8218;

architecture SYN_ARCHSTRUCT of mux21_8218 is

   component nd2_24652
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24653
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24654
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8218
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8218 port map( A => S, Y => n_S);
   NAND1 : nd2_24654 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24653 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24652 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8217 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8217;

architecture SYN_ARCHSTRUCT of mux21_8217 is

   component nd2_24649
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24650
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24651
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8217
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8217 port map( A => S, Y => n_S);
   NAND1 : nd2_24651 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24650 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24649 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8216 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8216;

architecture SYN_ARCHSTRUCT of mux21_8216 is

   component nd2_24646
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24647
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24648
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8216
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8216 port map( A => S, Y => n_S);
   NAND1 : nd2_24648 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24647 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24646 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8215 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8215;

architecture SYN_ARCHSTRUCT of mux21_8215 is

   component nd2_24643
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24644
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24645
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8215
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8215 port map( A => S, Y => n_S);
   NAND1 : nd2_24645 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24644 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24643 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8214 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8214;

architecture SYN_ARCHSTRUCT of mux21_8214 is

   component nd2_24640
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24641
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24642
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8214
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8214 port map( A => S, Y => n_S);
   NAND1 : nd2_24642 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24641 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24640 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8213 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8213;

architecture SYN_ARCHSTRUCT of mux21_8213 is

   component nd2_24637
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24638
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24639
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8213
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8213 port map( A => S, Y => n_S);
   NAND1 : nd2_24639 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24638 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24637 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8212 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8212;

architecture SYN_ARCHSTRUCT of mux21_8212 is

   component nd2_24634
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24635
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24636
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8212
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8212 port map( A => S, Y => n_S);
   NAND1 : nd2_24636 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24635 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24634 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8211 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8211;

architecture SYN_ARCHSTRUCT of mux21_8211 is

   component nd2_24631
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24632
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24633
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8211
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8211 port map( A => S, Y => n_S);
   NAND1 : nd2_24633 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24632 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24631 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8210 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8210;

architecture SYN_ARCHSTRUCT of mux21_8210 is

   component nd2_24628
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24629
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24630
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8210
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8210 port map( A => S, Y => n_S);
   NAND1 : nd2_24630 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24629 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24628 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8209 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8209;

architecture SYN_ARCHSTRUCT of mux21_8209 is

   component nd2_24625
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24626
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24627
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8209
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8209 port map( A => S, Y => n_S);
   NAND1 : nd2_24627 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24626 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24625 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8208 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8208;

architecture SYN_ARCHSTRUCT of mux21_8208 is

   component nd2_24622
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24623
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24624
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8208
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8208 port map( A => S, Y => n_S);
   NAND1 : nd2_24624 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24623 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24622 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8207 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8207;

architecture SYN_ARCHSTRUCT of mux21_8207 is

   component nd2_24619
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24620
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24621
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8207
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8207 port map( A => S, Y => n_S);
   NAND1 : nd2_24621 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24620 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24619 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8206 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8206;

architecture SYN_ARCHSTRUCT of mux21_8206 is

   component nd2_24616
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24617
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24618
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8206
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8206 port map( A => S, Y => n_S);
   NAND1 : nd2_24618 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24617 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24616 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8205 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8205;

architecture SYN_ARCHSTRUCT of mux21_8205 is

   component nd2_24613
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24614
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24615
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8205
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8205 port map( A => S, Y => n_S);
   NAND1 : nd2_24615 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24614 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24613 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8204 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8204;

architecture SYN_ARCHSTRUCT of mux21_8204 is

   component nd2_24610
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24611
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24612
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8204
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8204 port map( A => S, Y => n_S);
   NAND1 : nd2_24612 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24611 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24610 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8203 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8203;

architecture SYN_ARCHSTRUCT of mux21_8203 is

   component nd2_24607
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24608
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24609
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8203
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8203 port map( A => S, Y => n_S);
   NAND1 : nd2_24609 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24608 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24607 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8202 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8202;

architecture SYN_ARCHSTRUCT of mux21_8202 is

   component nd2_24604
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24605
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24606
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8202
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8202 port map( A => S, Y => n_S);
   NAND1 : nd2_24606 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24605 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24604 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8201 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8201;

architecture SYN_ARCHSTRUCT of mux21_8201 is

   component nd2_24601
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24602
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24603
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8201
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8201 port map( A => S, Y => n_S);
   NAND1 : nd2_24603 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24602 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24601 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8200 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8200;

architecture SYN_ARCHSTRUCT of mux21_8200 is

   component nd2_24598
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24599
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24600
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8200
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8200 port map( A => S, Y => n_S);
   NAND1 : nd2_24600 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24599 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24598 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8199 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8199;

architecture SYN_ARCHSTRUCT of mux21_8199 is

   component nd2_24595
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24596
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24597
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8199
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8199 port map( A => S, Y => n_S);
   NAND1 : nd2_24597 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24596 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24595 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8198 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8198;

architecture SYN_ARCHSTRUCT of mux21_8198 is

   component nd2_24592
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24593
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24594
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8198
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8198 port map( A => S, Y => n_S);
   NAND1 : nd2_24594 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24593 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24592 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8197 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8197;

architecture SYN_ARCHSTRUCT of mux21_8197 is

   component nd2_24589
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24590
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24591
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8197
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8197 port map( A => S, Y => n_S);
   NAND1 : nd2_24591 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24590 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24589 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8196 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8196;

architecture SYN_ARCHSTRUCT of mux21_8196 is

   component nd2_24586
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24587
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24588
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8196
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8196 port map( A => S, Y => n_S);
   NAND1 : nd2_24588 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24587 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24586 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8195 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8195;

architecture SYN_ARCHSTRUCT of mux21_8195 is

   component nd2_24583
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24584
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24585
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8195
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8195 port map( A => S, Y => n_S);
   NAND1 : nd2_24585 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24584 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24583 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8194 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8194;

architecture SYN_ARCHSTRUCT of mux21_8194 is

   component nd2_24580
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24581
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24582
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8194
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8194 port map( A => S, Y => n_S);
   NAND1 : nd2_24582 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24581 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24580 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8193 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8193;

architecture SYN_ARCHSTRUCT of mux21_8193 is

   component nd2_24577
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24578
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24579
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8193
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8193 port map( A => S, Y => n_S);
   NAND1 : nd2_24579 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24578 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24577 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8192 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8192;

architecture SYN_ARCHSTRUCT of mux21_8192 is

   component nd2_24574
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24575
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24576
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8192
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8192 port map( A => S, Y => n_S);
   NAND1 : nd2_24576 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24575 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24574 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8191 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8191;

architecture SYN_ARCHSTRUCT of mux21_8191 is

   component nd2_24571
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24572
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24573
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8191
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8191 port map( A => S, Y => n_S);
   NAND1 : nd2_24573 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24572 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24571 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8190 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8190;

architecture SYN_ARCHSTRUCT of mux21_8190 is

   component nd2_24568
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24569
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24570
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8190
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8190 port map( A => S, Y => n_S);
   NAND1 : nd2_24570 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24569 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24568 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8189 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8189;

architecture SYN_ARCHSTRUCT of mux21_8189 is

   component nd2_24565
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24566
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24567
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8189
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8189 port map( A => S, Y => n_S);
   NAND1 : nd2_24567 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24566 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24565 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8188 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8188;

architecture SYN_ARCHSTRUCT of mux21_8188 is

   component nd2_24562
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24563
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24564
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8188
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8188 port map( A => S, Y => n_S);
   NAND1 : nd2_24564 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24563 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24562 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8187 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8187;

architecture SYN_ARCHSTRUCT of mux21_8187 is

   component nd2_24559
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24560
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24561
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8187
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8187 port map( A => S, Y => n_S);
   NAND1 : nd2_24561 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24560 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24559 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8186 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8186;

architecture SYN_ARCHSTRUCT of mux21_8186 is

   component nd2_24556
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24557
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24558
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8186
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8186 port map( A => S, Y => n_S);
   NAND1 : nd2_24558 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24557 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24556 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8185 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8185;

architecture SYN_ARCHSTRUCT of mux21_8185 is

   component nd2_24553
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24554
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24555
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8185
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8185 port map( A => S, Y => n_S);
   NAND1 : nd2_24555 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24554 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24553 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8184 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8184;

architecture SYN_ARCHSTRUCT of mux21_8184 is

   component nd2_24550
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24551
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24552
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8184
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8184 port map( A => S, Y => n_S);
   NAND1 : nd2_24552 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24551 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24550 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8183 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8183;

architecture SYN_ARCHSTRUCT of mux21_8183 is

   component nd2_24547
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24548
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24549
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8183
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8183 port map( A => S, Y => n_S);
   NAND1 : nd2_24549 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24548 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24547 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8182 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8182;

architecture SYN_ARCHSTRUCT of mux21_8182 is

   component nd2_24544
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24545
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24546
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8182
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8182 port map( A => S, Y => n_S);
   NAND1 : nd2_24546 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24545 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24544 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8181 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8181;

architecture SYN_ARCHSTRUCT of mux21_8181 is

   component nd2_24541
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24542
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24543
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8181
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8181 port map( A => S, Y => n_S);
   NAND1 : nd2_24543 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24542 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24541 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8180 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8180;

architecture SYN_ARCHSTRUCT of mux21_8180 is

   component nd2_24538
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24539
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24540
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8180
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8180 port map( A => S, Y => n_S);
   NAND1 : nd2_24540 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24539 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24538 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8179 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8179;

architecture SYN_ARCHSTRUCT of mux21_8179 is

   component nd2_24535
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24536
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24537
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8179
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8179 port map( A => S, Y => n_S);
   NAND1 : nd2_24537 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24536 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24535 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8178 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8178;

architecture SYN_ARCHSTRUCT of mux21_8178 is

   component nd2_24532
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24533
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24534
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8178
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8178 port map( A => S, Y => n_S);
   NAND1 : nd2_24534 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24533 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24532 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8177 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8177;

architecture SYN_ARCHSTRUCT of mux21_8177 is

   component nd2_24529
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24530
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24531
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8177
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8177 port map( A => S, Y => n_S);
   NAND1 : nd2_24531 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24530 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24529 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8176 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8176;

architecture SYN_ARCHSTRUCT of mux21_8176 is

   component nd2_24526
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24527
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24528
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8176
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8176 port map( A => S, Y => n_S);
   NAND1 : nd2_24528 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24527 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24526 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8175 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8175;

architecture SYN_ARCHSTRUCT of mux21_8175 is

   component nd2_24523
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24524
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24525
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8175
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8175 port map( A => S, Y => n_S);
   NAND1 : nd2_24525 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24524 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24523 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8174 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8174;

architecture SYN_ARCHSTRUCT of mux21_8174 is

   component nd2_24520
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24521
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24522
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8174
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8174 port map( A => S, Y => n_S);
   NAND1 : nd2_24522 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24521 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24520 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8173 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8173;

architecture SYN_ARCHSTRUCT of mux21_8173 is

   component nd2_24517
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24518
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24519
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8173
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8173 port map( A => S, Y => n_S);
   NAND1 : nd2_24519 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24518 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24517 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8172 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8172;

architecture SYN_ARCHSTRUCT_architecture of mux21_8172 is

   component nd2_24514
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24515
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24516
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8172
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8172 port map( A => S, Y => n_S);
   NAND1 : nd2_24516 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24515 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24514 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8171 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8171;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8171 is

   component nd2_24511
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24512
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24513
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8171
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8171 port map( A => S, Y => n_S);
   NAND1 : nd2_24513 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24512 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24511 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8170 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8170;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8170 is

   component nd2_24508
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24509
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24510
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8170
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8170 port map( A => S, Y => n_S);
   NAND1 : nd2_24510 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24509 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24508 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8169 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8169;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8169 is

   component nd2_24505
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24506
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24507
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8169
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8169 port map( A => S, Y => n_S);
   NAND1 : nd2_24507 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24506 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24505 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8168 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8168;

architecture SYN_ARCHSTRUCT_architecture of mux21_8168 is

   component nd2_24502
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24503
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24504
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8168
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8168 port map( A => S, Y => n_S);
   NAND1 : nd2_24504 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24503 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24502 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8167 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8167;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8167 is

   component nd2_24499
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24500
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24501
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8167
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8167 port map( A => S, Y => n_S);
   NAND1 : nd2_24501 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24500 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24499 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8166 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8166;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8166 is

   component nd2_24496
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24497
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24498
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8166
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8166 port map( A => S, Y => n_S);
   NAND1 : nd2_24498 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24497 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24496 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8165 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8165;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8165 is

   component nd2_24493
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24494
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24495
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8165
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8165 port map( A => S, Y => n_S);
   NAND1 : nd2_24495 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24494 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24493 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8164 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8164;

architecture SYN_ARCHSTRUCT_architecture of mux21_8164 is

   component nd2_24490
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24491
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24492
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8164
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8164 port map( A => S, Y => n_S);
   NAND1 : nd2_24492 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24491 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24490 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8163 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8163;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8163 is

   component nd2_24487
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24488
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24489
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8163
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8163 port map( A => S, Y => n_S);
   NAND1 : nd2_24489 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24488 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24487 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8162 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8162;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8162 is

   component nd2_24484
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24485
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24486
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8162
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8162 port map( A => S, Y => n_S);
   NAND1 : nd2_24486 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24485 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24484 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8161 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8161;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8161 is

   component nd2_24481
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24482
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24483
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8161
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8161 port map( A => S, Y => n_S);
   NAND1 : nd2_24483 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24482 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24481 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8160 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8160;

architecture SYN_ARCHSTRUCT_architecture of mux21_8160 is

   component nd2_24478
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24479
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24480
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8160
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8160 port map( A => S, Y => n_S);
   NAND1 : nd2_24480 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24479 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24478 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8159 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8159;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8159 is

   component nd2_24475
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24476
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24477
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8159
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8159 port map( A => S, Y => n_S);
   NAND1 : nd2_24477 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24476 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24475 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8158 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8158;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8158 is

   component nd2_24472
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24473
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24474
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8158
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8158 port map( A => S, Y => n_S);
   NAND1 : nd2_24474 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24473 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24472 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8157 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8157;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8157 is

   component nd2_24469
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24470
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24471
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8157
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8157 port map( A => S, Y => n_S);
   NAND1 : nd2_24471 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24470 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24469 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8156 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8156;

architecture SYN_ARCHSTRUCT_architecture of mux21_8156 is

   component nd2_24466
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24467
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24468
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8156
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8156 port map( A => S, Y => n_S);
   NAND1 : nd2_24468 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24467 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24466 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8155 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8155;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8155 is

   component nd2_24463
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24464
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24465
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8155
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8155 port map( A => S, Y => n_S);
   NAND1 : nd2_24465 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24464 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24463 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8154 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8154;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8154 is

   component nd2_24460
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24461
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24462
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8154
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8154 port map( A => S, Y => n_S);
   NAND1 : nd2_24462 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24461 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24460 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8153 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8153;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8153 is

   component nd2_24457
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24458
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24459
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8153
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8153 port map( A => S, Y => n_S);
   NAND1 : nd2_24459 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24458 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24457 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8152 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8152;

architecture SYN_ARCHSTRUCT_architecture of mux21_8152 is

   component nd2_24454
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24455
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24456
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8152
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8152 port map( A => S, Y => n_S);
   NAND1 : nd2_24456 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24455 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24454 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8151 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8151;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8151 is

   component nd2_24451
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24452
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24453
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8151
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8151 port map( A => S, Y => n_S);
   NAND1 : nd2_24453 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24452 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24451 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8150 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8150;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8150 is

   component nd2_24448
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24449
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24450
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8150
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8150 port map( A => S, Y => n_S);
   NAND1 : nd2_24450 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24449 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24448 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8149 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8149;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8149 is

   component nd2_24445
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24446
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24447
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8149
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8149 port map( A => S, Y => n_S);
   NAND1 : nd2_24447 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24446 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24445 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8148 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8148;

architecture SYN_ARCHSTRUCT_architecture of mux21_8148 is

   component nd2_24442
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24443
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24444
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8148
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8148 port map( A => S, Y => n_S);
   NAND1 : nd2_24444 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24443 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24442 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8147 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8147;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8147 is

   component nd2_24439
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24440
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24441
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8147
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8147 port map( A => S, Y => n_S);
   NAND1 : nd2_24441 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24440 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24439 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8146 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8146;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8146 is

   component nd2_24436
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24437
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24438
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8146
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8146 port map( A => S, Y => n_S);
   NAND1 : nd2_24438 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24437 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24436 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8145 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8145;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8145 is

   component nd2_24433
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24434
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24435
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8145
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8145 port map( A => S, Y => n_S);
   NAND1 : nd2_24435 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24434 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24433 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8144 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8144;

architecture SYN_ARCHSTRUCT_architecture of mux21_8144 is

   component nd2_24430
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24431
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24432
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8144
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8144 port map( A => S, Y => n_S);
   NAND1 : nd2_24432 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24431 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24430 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8143 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8143;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8143 is

   component nd2_24427
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24428
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24429
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8143
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8143 port map( A => S, Y => n_S);
   NAND1 : nd2_24429 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24428 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24427 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8142 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8142;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8142 is

   component nd2_24424
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24425
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24426
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8142
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8142 port map( A => S, Y => n_S);
   NAND1 : nd2_24426 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24425 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24424 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8141 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8141;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8141 is

   component nd2_24421
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24422
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24423
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8141
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8141 port map( A => S, Y => n_S);
   NAND1 : nd2_24423 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24422 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24421 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8140 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8140;

architecture SYN_ARCHSTRUCT_architecture of mux21_8140 is

   component nd2_24418
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24419
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24420
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8140
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8140 port map( A => S, Y => n_S);
   NAND1 : nd2_24420 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24419 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24418 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8139 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8139;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8139 is

   component nd2_24415
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24416
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24417
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8139
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8139 port map( A => S, Y => n_S);
   NAND1 : nd2_24417 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24416 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24415 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8138 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8138;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8138 is

   component nd2_24412
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24413
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24414
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8138
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8138 port map( A => S, Y => n_S);
   NAND1 : nd2_24414 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24413 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24412 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8137 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8137;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8137 is

   component nd2_24409
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24410
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24411
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8137
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8137 port map( A => S, Y => n_S);
   NAND1 : nd2_24411 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24410 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24409 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8136 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8136;

architecture SYN_ARCHSTRUCT_architecture of mux21_8136 is

   component nd2_24406
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24407
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24408
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8136
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8136 port map( A => S, Y => n_S);
   NAND1 : nd2_24408 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24407 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24406 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8135 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8135;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8135 is

   component nd2_24403
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24404
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24405
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8135
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8135 port map( A => S, Y => n_S);
   NAND1 : nd2_24405 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24404 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24403 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8134 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8134;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8134 is

   component nd2_24400
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24401
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24402
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8134
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8134 port map( A => S, Y => n_S);
   NAND1 : nd2_24402 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24401 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24400 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8133 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8133;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8133 is

   component nd2_24397
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24398
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24399
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8133
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8133 port map( A => S, Y => n_S);
   NAND1 : nd2_24399 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24398 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24397 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8132 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8132;

architecture SYN_ARCHSTRUCT_architecture of mux21_8132 is

   component nd2_24394
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24395
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24396
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8132
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8132 port map( A => S, Y => n_S);
   NAND1 : nd2_24396 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24395 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24394 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8131 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8131;

architecture SYN_ARCHSTRUCT_architecture2 of mux21_8131 is

   component nd2_24391
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24392
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24393
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8131
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8131 port map( A => S, Y => n_S);
   NAND1 : nd2_24393 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24392 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24391 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8130 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8130;

architecture SYN_ARCHSTRUCT_architecture3 of mux21_8130 is

   component nd2_24388
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24389
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24390
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8130
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8130 port map( A => S, Y => n_S);
   NAND1 : nd2_24390 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24389 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24388 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8129 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8129;

architecture SYN_ARCHSTRUCT_architecture4 of mux21_8129 is

   component nd2_24385
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24386
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24387
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8129
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2 : std_logic;

begin
   
   NOT1 : iv_8129 port map( A => S, Y => n_S);
   NAND1 : nd2_24387 port map( A => A, B => S, Y => s1);
   NAND2 : nd2_24386 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_24385 port map( A => s1, B => s2, Y => Y);

end SYN_ARCHSTRUCT_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity sum_generator_N16_Nbit_blocks4_2 is

   port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  Carry 
         : in std_logic_vector (3 downto 0);  S : out std_logic_vector (15 
         downto 0);  Cout : out std_logic);

end sum_generator_N16_Nbit_blocks4_2;

architecture SYN_ARCHSTRUCT of sum_generator_N16_Nbit_blocks4_2 is

   component carry_select_block_N4_245
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_246
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_247
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_248
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   Cout <= Carry(3);
   
   CSB_1 : carry_select_block_N4_248 port map( Cin => Cin, A(3) => A(3), A(2) 
                           => A(2), A(1) => A(1), A(0) => A(0), B(3) => B(3), 
                           B(2) => B(2), B(1) => B(1), B(0) => B(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSB_2 : carry_select_block_N4_247 port map( Cin => Carry(0), A(3) => A(7), 
                           A(2) => A(6), A(1) => A(5), A(0) => A(4), B(3) => 
                           B(7), B(2) => B(6), B(1) => B(5), B(0) => B(4), S(3)
                           => S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CSB_3 : carry_select_block_N4_246 port map( Cin => Carry(1), A(3) => A(11), 
                           A(2) => A(10), A(1) => A(9), A(0) => A(8), B(3) => 
                           B(11), B(2) => B(10), B(1) => B(9), B(0) => B(8), 
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   CSB_4 : carry_select_block_N4_245 port map( Cin => Carry(2), A(3) => A(15), 
                           A(2) => A(14), A(1) => A(13), A(0) => A(12), B(3) =>
                           B(15), B(2) => B(14), B(1) => B(13), B(0) => B(12), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity sum_generator_N16_Nbit_blocks4_1 is

   port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  Carry 
         : in std_logic_vector (3 downto 0);  S : out std_logic_vector (15 
         downto 0);  Cout : out std_logic);

end sum_generator_N16_Nbit_blocks4_1;

architecture SYN_ARCHSTRUCT of sum_generator_N16_Nbit_blocks4_1 is

   component carry_select_block_N4_241
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_242
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_243
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_244
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   Cout <= Carry(3);
   
   CSB_1 : carry_select_block_N4_244 port map( Cin => Cin, A(3) => A(3), A(2) 
                           => A(2), A(1) => A(1), A(0) => A(0), B(3) => B(3), 
                           B(2) => B(2), B(1) => B(1), B(0) => B(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSB_2 : carry_select_block_N4_243 port map( Cin => Carry(0), A(3) => A(7), 
                           A(2) => A(6), A(1) => A(5), A(0) => A(4), B(3) => 
                           B(7), B(2) => B(6), B(1) => B(5), B(0) => B(4), S(3)
                           => S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CSB_3 : carry_select_block_N4_242 port map( Cin => Carry(1), A(3) => A(11), 
                           A(2) => A(10), A(1) => A(9), A(0) => A(8), B(3) => 
                           B(11), B(2) => B(10), B(1) => B(9), B(0) => B(8), 
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   CSB_4 : carry_select_block_N4_241 port map( Cin => Carry(2), A(3) => A(15), 
                           A(2) => A(14), A(1) => A(13), A(0) => A(12), B(3) =>
                           B(15), B(2) => B(14), B(1) => B(13), B(0) => B(12), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_generator_N16_carry_range4_2 is

   port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C : 
         out std_logic_vector (4 downto 0));

end carry_generator_N16_carry_range4_2;

architecture SYN_ARCHSTRUCT of carry_generator_N16_carry_range4_2 is

   component carry_generator_sparse_tree_N16_carry_range4_2
      port( P, G : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C :
            out std_logic_vector (4 downto 0));
   end component;
   
   component pg_network_N16_2
      port( A, B : in std_logic_vector (15 downto 0);  P, G : out 
            std_logic_vector (15 downto 0));
   end component;
   
   signal P_15_port, P_14_port, P_13_port, P_12_port, P_11_port, P_10_port, 
      P_9_port, P_8_port, P_7_port, P_6_port, P_5_port, P_4_port, P_3_port, 
      P_2_port, P_1_port, P_0_port, G_15_port, G_14_port, G_13_port, G_12_port,
      G_11_port, G_10_port, G_9_port, G_8_port, G_7_port, G_6_port, G_5_port, 
      G_4_port, G_3_port, G_2_port, G_1_port, G_0_port : std_logic;

begin
   
   PG_NET : pg_network_N16_2 port map( A(15) => A(15), A(14) => A(14), A(13) =>
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), P(15) => P_15_port
                           , P(14) => P_14_port, P(13) => P_13_port, P(12) => 
                           P_12_port, P(11) => P_11_port, P(10) => P_10_port, 
                           P(9) => P_9_port, P(8) => P_8_port, P(7) => P_7_port
                           , P(6) => P_6_port, P(5) => P_5_port, P(4) => 
                           P_4_port, P(3) => P_3_port, P(2) => P_2_port, P(1) 
                           => P_1_port, P(0) => P_0_port, G(15) => G_15_port, 
                           G(14) => G_14_port, G(13) => G_13_port, G(12) => 
                           G_12_port, G(11) => G_11_port, G(10) => G_10_port, 
                           G(9) => G_9_port, G(8) => G_8_port, G(7) => G_7_port
                           , G(6) => G_6_port, G(5) => G_5_port, G(4) => 
                           G_4_port, G(3) => G_3_port, G(2) => G_2_port, G(1) 
                           => G_1_port, G(0) => G_0_port);
   CG : carry_generator_sparse_tree_N16_carry_range4_2 port map( P(15) => 
                           P_15_port, P(14) => P_14_port, P(13) => P_13_port, 
                           P(12) => P_12_port, P(11) => P_11_port, P(10) => 
                           P_10_port, P(9) => P_9_port, P(8) => P_8_port, P(7) 
                           => P_7_port, P(6) => P_6_port, P(5) => P_5_port, 
                           P(4) => P_4_port, P(3) => P_3_port, P(2) => P_2_port
                           , P(1) => P_1_port, P(0) => P_0_port, G(15) => 
                           G_15_port, G(14) => G_14_port, G(13) => G_13_port, 
                           G(12) => G_12_port, G(11) => G_11_port, G(10) => 
                           G_10_port, G(9) => G_9_port, G(8) => G_8_port, G(7) 
                           => G_7_port, G(6) => G_6_port, G(5) => G_5_port, 
                           G(4) => G_4_port, G(3) => G_3_port, G(2) => G_2_port
                           , G(1) => G_1_port, G(0) => G_0_port, Cin => Cin, 
                           C(4) => C(4), C(3) => C(3), C(2) => C(2), C(1) => 
                           C(1), C(0) => C(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_generator_N16_carry_range4_1 is

   port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C : 
         out std_logic_vector (4 downto 0));

end carry_generator_N16_carry_range4_1;

architecture SYN_ARCHSTRUCT of carry_generator_N16_carry_range4_1 is

   component carry_generator_sparse_tree_N16_carry_range4_1
      port( P, G : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C :
            out std_logic_vector (4 downto 0));
   end component;
   
   component pg_network_N16_1
      port( A, B : in std_logic_vector (15 downto 0);  P, G : out 
            std_logic_vector (15 downto 0));
   end component;
   
   signal P_15_port, P_14_port, P_13_port, P_12_port, P_11_port, P_10_port, 
      P_9_port, P_8_port, P_7_port, P_6_port, P_5_port, P_4_port, P_3_port, 
      P_2_port, P_1_port, P_0_port, G_15_port, G_14_port, G_13_port, G_12_port,
      G_11_port, G_10_port, G_9_port, G_8_port, G_7_port, G_6_port, G_5_port, 
      G_4_port, G_3_port, G_2_port, G_1_port, G_0_port : std_logic;

begin
   
   PG_NET : pg_network_N16_1 port map( A(15) => A(15), A(14) => A(14), A(13) =>
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), P(15) => P_15_port
                           , P(14) => P_14_port, P(13) => P_13_port, P(12) => 
                           P_12_port, P(11) => P_11_port, P(10) => P_10_port, 
                           P(9) => P_9_port, P(8) => P_8_port, P(7) => P_7_port
                           , P(6) => P_6_port, P(5) => P_5_port, P(4) => 
                           P_4_port, P(3) => P_3_port, P(2) => P_2_port, P(1) 
                           => P_1_port, P(0) => P_0_port, G(15) => G_15_port, 
                           G(14) => G_14_port, G(13) => G_13_port, G(12) => 
                           G_12_port, G(11) => G_11_port, G(10) => G_10_port, 
                           G(9) => G_9_port, G(8) => G_8_port, G(7) => G_7_port
                           , G(6) => G_6_port, G(5) => G_5_port, G(4) => 
                           G_4_port, G(3) => G_3_port, G(2) => G_2_port, G(1) 
                           => G_1_port, G(0) => G_0_port);
   CG : carry_generator_sparse_tree_N16_carry_range4_1 port map( P(15) => 
                           P_15_port, P(14) => P_14_port, P(13) => P_13_port, 
                           P(12) => P_12_port, P(11) => P_11_port, P(10) => 
                           P_10_port, P(9) => P_9_port, P(8) => P_8_port, P(7) 
                           => P_7_port, P(6) => P_6_port, P(5) => P_5_port, 
                           P(4) => P_4_port, P(3) => P_3_port, P(2) => P_2_port
                           , P(1) => P_1_port, P(0) => P_0_port, G(15) => 
                           G_15_port, G(14) => G_14_port, G(13) => G_13_port, 
                           G(12) => G_12_port, G(11) => G_11_port, G(10) => 
                           G_10_port, G(9) => G_9_port, G(8) => G_8_port, G(7) 
                           => G_7_port, G(6) => G_6_port, G(5) => G_5_port, 
                           G(4) => G_4_port, G(3) => G_3_port, G(2) => G_2_port
                           , G(1) => G_1_port, G(0) => G_0_port, Cin => Cin, 
                           C(4) => C(4), C(3) => C(3), C(2) => C(2), C(1) => 
                           C(1), C(0) => C(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_27 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_27;

architecture SYN_ARCHSTRUCT of muxN1_N16_27 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8593
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8594
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8595
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8596
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8597
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8598
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8599
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8600
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8601
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8602
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8603
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8604
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8605
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8606
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8607
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8608
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8608 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8607 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8606 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8605 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8604 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8603 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8602 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8601 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8600 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8599 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8598 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8597 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8596 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8595 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8594 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8593 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n2);
   U2 : BUF_X1 port map( A => n1, Z => n3);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_26 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_26;

architecture SYN_ARCHSTRUCT of muxN1_N16_26 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8577
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8578
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8579
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8580
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8581
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8582
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8583
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8584
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8585
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8586
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8587
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8588
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8589
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8590
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8591
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8592
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8592 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8591 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8590 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8589 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8588 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8587 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8586 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8585 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8584 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8583 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8582 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8581 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8580 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8579 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8578 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8577 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n2);
   U2 : BUF_X1 port map( A => n1, Z => n3);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_25 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_25;

architecture SYN_ARCHSTRUCT of muxN1_N16_25 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8561
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8562
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8563
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8564
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8565
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8566
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8567
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8568
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8569
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8570
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8571
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8572
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8573
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8574
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8575
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8576
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8576 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8575 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8574 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8573 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8572 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8571 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8570 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8569 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8568 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8567 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8566 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8565 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8564 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8563 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8562 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8561 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n2);
   U2 : BUF_X1 port map( A => n1, Z => n3);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_24 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_24;

architecture SYN_ARCHSTRUCT of muxN1_N16_24 is

   component mux21_8545
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8546
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8547
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8548
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8549
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8550
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8551
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8552
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8553
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8554
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8555
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8556
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8557
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8558
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8559
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8560
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8560 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8559 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8558 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8557 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8556 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8555 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8554 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8553 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8552 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8551 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8550 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8549 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8548 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8547 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8546 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8545 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_23 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_23;

architecture SYN_ARCHSTRUCT of muxN1_N16_23 is

   component mux21_8529
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8530
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8531
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8532
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8533
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8534
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8535
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8536
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8537
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8538
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8539
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8540
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8541
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8542
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8543
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8544
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8544 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8543 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8542 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8541 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8540 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8539 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8538 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8537 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8536 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8535 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8534 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8533 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8532 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8531 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8530 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8529 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_22 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_22;

architecture SYN_ARCHSTRUCT of muxN1_N16_22 is

   component mux21_8513
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8514
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8515
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8516
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8517
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8518
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8519
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8520
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8521
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8522
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8523
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8524
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8525
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8526
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8527
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8528
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8528 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8527 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8526 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8525 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8524 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8523 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8522 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8521 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8520 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8519 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8518 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8517 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8516 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8515 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8514 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8513 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_21 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_21;

architecture SYN_ARCHSTRUCT of muxN1_N16_21 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8497
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8498
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8499
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8500
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8501
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8502
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8503
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8504
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8505
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8506
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8507
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8508
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8509
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8510
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8511
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8512
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8512 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8511 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8510 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8509 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8508 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8507 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8506 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8505 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8504 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8503 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8502 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8501 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8500 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8499 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8498 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8497 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_20 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_20;

architecture SYN_ARCHSTRUCT of muxN1_N16_20 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8481
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8482
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8483
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8484
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8485
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8486
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8487
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8488
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8489
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8490
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8491
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8492
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8493
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8494
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8495
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8496
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8496 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8495 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8494 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8493 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8492 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8491 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8490 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8489 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8488 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8487 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8486 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8485 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8484 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8483 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8482 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8481 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_19 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_19;

architecture SYN_ARCHSTRUCT of muxN1_N16_19 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8465
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8466
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8467
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8468
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8469
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8470
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8471
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8472
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8473
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8474
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8475
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8476
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8477
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8478
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8479
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8480
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8480 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8479 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8478 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8477 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8476 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8475 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8474 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8473 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8472 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8471 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8470 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8469 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8468 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8467 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8466 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8465 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_18 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_18;

architecture SYN_ARCHSTRUCT of muxN1_N16_18 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8449
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8450
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8451
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8452
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8453
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8454
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8455
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8456
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8457
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8458
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8459
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8460
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8461
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8462
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8463
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8464
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8464 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8463 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8462 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8461 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8460 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8459 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8458 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8457 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8456 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8455 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8454 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8453 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8452 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8451 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8450 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8449 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_17 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_17;

architecture SYN_ARCHSTRUCT of muxN1_N16_17 is

   component mux21_8433
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8434
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8435
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8436
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8437
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8438
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8439
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8440
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8441
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8442
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8443
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8444
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8445
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8446
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8447
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8448
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8448 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8447 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8446 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8445 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8444 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8443 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8442 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8441 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8440 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8439 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8438 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8437 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8436 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8435 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8434 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8433 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_16 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_16;

architecture SYN_ARCHSTRUCT of muxN1_N16_16 is

   component mux21_8417
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8418
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8419
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8420
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8421
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8422
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8423
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8424
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8425
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8426
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8427
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8428
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8429
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8430
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8431
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8432
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8432 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8431 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8430 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8429 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8428 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8427 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8426 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8425 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8424 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8423 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8422 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8421 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8420 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8419 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8418 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8417 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_15 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_15;

architecture SYN_ARCHSTRUCT of muxN1_N16_15 is

   component mux21_8401
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8402
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8403
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8404
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8405
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8406
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8407
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8408
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8409
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8410
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8411
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8412
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8413
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8414
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8415
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8416
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8416 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8415 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8414 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8413 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8412 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8411 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8410 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8409 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8408 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8407 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8406 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8405 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8404 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8403 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8402 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8401 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_14 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_14;

architecture SYN_ARCHSTRUCT of muxN1_N16_14 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8385
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8386
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8387
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8388
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8389
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8390
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8391
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8392
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8393
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8394
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8395
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8396
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8397
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8398
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8399
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8400
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8400 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8399 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8398 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8397 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8396 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8395 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8394 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8393 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8392 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8391 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8390 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8389 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8388 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8387 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8386 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8385 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_13 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_13;

architecture SYN_ARCHSTRUCT of muxN1_N16_13 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8369
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8370
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8371
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8372
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8373
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8374
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8375
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8376
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8377
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8378
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8379
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8380
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8381
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8382
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8383
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8384
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8384 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8383 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8382 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8381 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8380 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8379 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8378 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8377 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8376 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8375 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8374 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8373 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8372 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8371 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8370 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8369 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_12 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_12;

architecture SYN_ARCHSTRUCT of muxN1_N16_12 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8353
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8354
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8355
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8356
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8357
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8358
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8359
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8360
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8361
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8362
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8363
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8364
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8365
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8366
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8367
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8368
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8368 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8367 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8366 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8365 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8364 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8363 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8362 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8361 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8360 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8359 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8358 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8357 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8356 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8355 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8354 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8353 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_11 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_11;

architecture SYN_ARCHSTRUCT of muxN1_N16_11 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8337
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8338
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8339
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8340
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8341
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8342
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8343
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8344
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8345
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8346
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8347
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8348
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8349
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8350
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8351
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8352
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8352 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8351 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8350 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8349 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8348 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8347 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8346 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8345 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8344 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8343 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8342 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8341 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8340 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8339 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8338 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8337 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_10 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_10;

architecture SYN_ARCHSTRUCT of muxN1_N16_10 is

   component mux21_8321
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8322
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8323
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8324
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8325
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8326
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8327
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8328
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8329
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8330
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8331
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8332
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8333
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8334
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8335
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8336
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8336 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8335 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8334 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8333 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8332 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8331 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8330 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8329 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8328 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8327 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8326 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8325 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8324 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8323 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8322 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8321 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_9 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_9;

architecture SYN_ARCHSTRUCT of muxN1_N16_9 is

   component mux21_8305
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8306
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8307
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8308
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8309
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8310
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8311
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8312
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8313
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8314
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8315
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8316
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8317
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8318
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8319
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8320
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8320 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8319 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8318 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8317 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8316 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8315 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8314 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8313 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8312 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8311 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8310 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8309 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8308 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8307 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8306 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8305 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_8 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_8;

architecture SYN_ARCHSTRUCT of muxN1_N16_8 is

   component mux21_8289
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8290
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8291
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8292
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8293
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8294
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8295
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8296
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8297
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8298
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8299
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8300
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8301
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8302
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8303
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8304
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8304 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8303 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8302 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8301 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8300 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8299 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8298 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8297 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8296 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8295 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8294 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8293 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8292 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8291 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8290 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8289 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_7 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_7;

architecture SYN_ARCHSTRUCT of muxN1_N16_7 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8273
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8274
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8275
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8276
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8277
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8278
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8279
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8280
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8281
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8282
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8283
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8284
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8285
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8286
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8287
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8288
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8288 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8287 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8286 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8285 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8284 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8283 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8282 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8281 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8280 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8279 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8278 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8277 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8276 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8275 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8274 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8273 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_6 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_6;

architecture SYN_ARCHSTRUCT of muxN1_N16_6 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8257
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8258
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8259
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8260
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8261
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8262
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8263
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8264
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8265
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8266
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8267
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8268
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8269
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8270
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8271
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8272
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8272 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8271 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8270 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8269 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8268 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8267 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8266 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8265 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8264 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8263 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8262 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8261 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8260 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8259 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8258 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8257 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_5 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_5;

architecture SYN_ARCHSTRUCT of muxN1_N16_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8241
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8242
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8243
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8244
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8245
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8246
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8247
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8248
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8249
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8250
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8251
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8252
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8253
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8254
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8255
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8256
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8256 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8255 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8254 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8253 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8252 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8251 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8250 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8249 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8248 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8247 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8246 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8245 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8244 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8243 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8242 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8241 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_4 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_4;

architecture SYN_ARCHSTRUCT of muxN1_N16_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8225
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8226
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8227
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8228
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8229
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8230
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8231
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8232
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8233
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8234
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8235
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8236
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8237
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8238
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8239
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8240
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8240 port map( A => A(0), B => B(0), S => n2, Y => Y(0));
   mux21_g_1 : mux21_8239 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8238 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8237 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8236 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8235 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8234 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8233 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8232 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8231 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8230 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8229 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8228 port map( A => A(12), B => B(12), S => n3, Y => 
                           Y(12));
   mux21_g_13 : mux21_8227 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8226 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8225 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n3);
   U2 : BUF_X1 port map( A => n1, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_3 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_3;

architecture SYN_ARCHSTRUCT of muxN1_N16_3 is

   component mux21_8209
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8210
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8211
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8212
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8213
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8214
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8215
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8216
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8217
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8218
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8219
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8220
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8221
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8222
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8223
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8224
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8224 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8223 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8222 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8221 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8220 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8219 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8218 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8217 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8216 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8215 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8214 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8213 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8212 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8211 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8210 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8209 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_2 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_2;

architecture SYN_ARCHSTRUCT of muxN1_N16_2 is

   component mux21_8193
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8194
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8195
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8196
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8197
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8198
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8199
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8200
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8201
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8202
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8203
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8204
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8205
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8206
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8207
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8208
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8208 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8207 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8206 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8205 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8204 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8203 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8202 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8201 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8200 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8199 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8198 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8197 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8196 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8195 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8194 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8193 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_1 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_1;

architecture SYN_ARCHSTRUCT of muxN1_N16_1 is

   component mux21_8177
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8178
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8179
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8180
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8181
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8182
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8183
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8184
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8185
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8186
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8187
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8188
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8189
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8190
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8191
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8192
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8192 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8191 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8190 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8189 port map( A => A(3), B => B(3), S => S, Y => Y(3));
   mux21_g_4 : mux21_8188 port map( A => A(4), B => B(4), S => S, Y => Y(4));
   mux21_g_5 : mux21_8187 port map( A => A(5), B => B(5), S => S, Y => Y(5));
   mux21_g_6 : mux21_8186 port map( A => A(6), B => B(6), S => S, Y => Y(6));
   mux21_g_7 : mux21_8185 port map( A => A(7), B => B(7), S => S, Y => Y(7));
   mux21_g_8 : mux21_8184 port map( A => A(8), B => B(8), S => S, Y => Y(8));
   mux21_g_9 : mux21_8183 port map( A => A(9), B => B(9), S => S, Y => Y(9));
   mux21_g_10 : mux21_8182 port map( A => A(10), B => B(10), S => S, Y => Y(10)
                           );
   mux21_g_11 : mux21_8181 port map( A => A(11), B => B(11), S => S, Y => Y(11)
                           );
   mux21_g_12 : mux21_8180 port map( A => A(12), B => B(12), S => S, Y => Y(12)
                           );
   mux21_g_13 : mux21_8179 port map( A => A(13), B => B(13), S => S, Y => Y(13)
                           );
   mux21_g_14 : mux21_8178 port map( A => A(14), B => B(14), S => S, Y => Y(14)
                           );
   mux21_g_15 : mux21_8177 port map( A => A(15), B => B(15), S => S, Y => Y(15)
                           );

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity booth_encoder_block_19 is

   port( Bi : in std_logic_vector (2 downto 0);  So : out std_logic_vector (2 
         downto 0));

end booth_encoder_block_19;

architecture SYN_DATAFLOW of booth_encoder_block_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U3 : INV_X4 port map( A => Bi(1), ZN => So(1));
   U4 : INV_X2 port map( A => Bi(2), ZN => So(2));
   U5 : INV_X1 port map( A => Bi(0), ZN => So(0));

end SYN_DATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity booth_encoder_block_18 is

   port( Bi : in std_logic_vector (2 downto 0);  So : out std_logic_vector (2 
         downto 0));

end booth_encoder_block_18;

architecture SYN_DATAFLOW of booth_encoder_block_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U3 : INV_X4 port map( A => Bi(1), ZN => So(1));
   U4 : INV_X2 port map( A => Bi(2), ZN => So(2));
   U5 : INV_X1 port map( A => Bi(0), ZN => So(0));

end SYN_DATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity booth_encoder_block_17 is

   port( Bi : in std_logic_vector (2 downto 0);  So : out std_logic_vector (2 
         downto 0));

end booth_encoder_block_17;

architecture SYN_DATAFLOW of booth_encoder_block_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U3 : INV_X4 port map( A => Bi(1), ZN => So(1));
   U4 : INV_X2 port map( A => Bi(2), ZN => So(2));
   U5 : INV_X1 port map( A => Bi(0), ZN => So(0));

end SYN_DATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity P4_adder_N16_Nbit_blocks4_2 is

   port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (15 downto 0);  Cout : out std_logic);

end P4_adder_N16_Nbit_blocks4_2;

architecture SYN_STRUCT of P4_adder_N16_Nbit_blocks4_2 is

   component sum_generator_N16_Nbit_blocks4_2
      port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  
            Carry : in std_logic_vector (3 downto 0);  S : out std_logic_vector
            (15 downto 0);  Cout : out std_logic);
   end component;
   
   component carry_generator_N16_carry_range4_2
      port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C :
            out std_logic_vector (4 downto 0));
   end component;
   
   signal Carries_4_port, Carries_3_port, Carries_2_port, Carries_1_port, 
      n_1118 : std_logic;

begin
   
   CG : carry_generator_N16_carry_range4_2 port map( A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), Cin 
                           => Cin, C(4) => Carries_4_port, C(3) => 
                           Carries_3_port, C(2) => Carries_2_port, C(1) => 
                           Carries_1_port, C(0) => n_1118);
   SG : sum_generator_N16_Nbit_blocks4_2 port map( A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), Cin 
                           => Cin, Carry(3) => Carries_4_port, Carry(2) => 
                           Carries_3_port, Carry(1) => Carries_2_port, Carry(0)
                           => Carries_1_port, S(15) => S(15), S(14) => S(14), 
                           S(13) => S(13), S(12) => S(12), S(11) => S(11), 
                           S(10) => S(10), S(9) => S(9), S(8) => S(8), S(7) => 
                           S(7), S(6) => S(6), S(5) => S(5), S(4) => S(4), S(3)
                           => S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0), 
                           Cout => Cout);

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity P4_adder_N16_Nbit_blocks4_1 is

   port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (15 downto 0);  Cout : out std_logic);

end P4_adder_N16_Nbit_blocks4_1;

architecture SYN_STRUCT of P4_adder_N16_Nbit_blocks4_1 is

   component sum_generator_N16_Nbit_blocks4_1
      port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  
            Carry : in std_logic_vector (3 downto 0);  S : out std_logic_vector
            (15 downto 0);  Cout : out std_logic);
   end component;
   
   component carry_generator_N16_carry_range4_1
      port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C :
            out std_logic_vector (4 downto 0));
   end component;
   
   signal Carries_4_port, Carries_3_port, Carries_2_port, Carries_1_port, 
      n_1119 : std_logic;

begin
   
   CG : carry_generator_N16_carry_range4_1 port map( A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), Cin 
                           => Cin, C(4) => Carries_4_port, C(3) => 
                           Carries_3_port, C(2) => Carries_2_port, C(1) => 
                           Carries_1_port, C(0) => n_1119);
   SG : sum_generator_N16_Nbit_blocks4_1 port map( A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), Cin 
                           => Cin, Carry(3) => Carries_4_port, Carry(2) => 
                           Carries_3_port, Carry(1) => Carries_2_port, Carry(0)
                           => Carries_1_port, S(15) => S(15), S(14) => S(14), 
                           S(13) => S(13), S(12) => S(12), S(11) => S(11), 
                           S(10) => S(10), S(9) => S(9), S(8) => S(8), S(7) => 
                           S(7), S(6) => S(6), S(5) => S(5), S(4) => S(4), S(3)
                           => S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0), 
                           Cout => Cout);

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux_8to1_N16_3 is

   port( A1, A2, A3, A4, A5, A6, A7, A8 : in std_logic_vector (15 downto 0);  S
         : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end mux_8to1_N16_3;

architecture SYN_ARCHSTRUCT of mux_8to1_N16_3 is

   component muxN1_N16_15
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_16
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_17
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_18
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_19
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_20
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_21
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   signal out1_15_port, out1_14_port, out1_13_port, out1_12_port, out1_11_port,
      out1_10_port, out1_9_port, out1_8_port, out1_7_port, out1_6_port, 
      out1_5_port, out1_4_port, out1_3_port, out1_2_port, out1_1_port, 
      out1_0_port, out2_15_port, out2_14_port, out2_13_port, out2_12_port, 
      out2_11_port, out2_10_port, out2_9_port, out2_8_port, out2_7_port, 
      out2_6_port, out2_5_port, out2_4_port, out2_3_port, out2_2_port, 
      out2_1_port, out2_0_port, out3_15_port, out3_14_port, out3_13_port, 
      out3_12_port, out3_11_port, out3_10_port, out3_9_port, out3_8_port, 
      out3_7_port, out3_6_port, out3_5_port, out3_4_port, out3_3_port, 
      out3_2_port, out3_1_port, out3_0_port, out4_15_port, out4_14_port, 
      out4_13_port, out4_12_port, out4_11_port, out4_10_port, out4_9_port, 
      out4_8_port, out4_7_port, out4_6_port, out4_5_port, out4_4_port, 
      out4_3_port, out4_2_port, out4_1_port, out4_0_port, out5_15_port, 
      out5_14_port, out5_13_port, out5_12_port, out5_11_port, out5_10_port, 
      out5_9_port, out5_8_port, out5_7_port, out5_6_port, out5_5_port, 
      out5_4_port, out5_3_port, out5_2_port, out5_1_port, out5_0_port, 
      out6_15_port, out6_14_port, out6_13_port, out6_12_port, out6_11_port, 
      out6_10_port, out6_9_port, out6_8_port, out6_7_port, out6_6_port, 
      out6_5_port, out6_4_port, out6_3_port, out6_2_port, out6_1_port, 
      out6_0_port : std_logic;

begin
   
   MUX1 : muxN1_N16_21 port map( A(15) => A1(15), A(14) => A1(14), A(13) => 
                           A1(13), A(12) => A1(12), A(11) => A1(11), A(10) => 
                           A1(10), A(9) => A1(9), A(8) => A1(8), A(7) => A1(7),
                           A(6) => A1(6), A(5) => A1(5), A(4) => A1(4), A(3) =>
                           A1(3), A(2) => A1(2), A(1) => A1(1), A(0) => A1(0), 
                           B(15) => A2(15), B(14) => A2(14), B(13) => A2(13), 
                           B(12) => A2(12), B(11) => A2(11), B(10) => A2(10), 
                           B(9) => A2(9), B(8) => A2(8), B(7) => A2(7), B(6) =>
                           A2(6), B(5) => A2(5), B(4) => A2(4), B(3) => A2(3), 
                           B(2) => A2(2), B(1) => A2(1), B(0) => A2(0), S => 
                           S(0), Y(15) => out1_15_port, Y(14) => out1_14_port, 
                           Y(13) => out1_13_port, Y(12) => out1_12_port, Y(11) 
                           => out1_11_port, Y(10) => out1_10_port, Y(9) => 
                           out1_9_port, Y(8) => out1_8_port, Y(7) => 
                           out1_7_port, Y(6) => out1_6_port, Y(5) => 
                           out1_5_port, Y(4) => out1_4_port, Y(3) => 
                           out1_3_port, Y(2) => out1_2_port, Y(1) => 
                           out1_1_port, Y(0) => out1_0_port);
   MUX2 : muxN1_N16_20 port map( A(15) => A3(15), A(14) => A3(14), A(13) => 
                           A3(13), A(12) => A3(12), A(11) => A3(11), A(10) => 
                           A3(10), A(9) => A3(9), A(8) => A3(8), A(7) => A3(7),
                           A(6) => A3(6), A(5) => A3(5), A(4) => A3(4), A(3) =>
                           A3(3), A(2) => A3(2), A(1) => A3(1), A(0) => A3(0), 
                           B(15) => A4(15), B(14) => A4(14), B(13) => A4(13), 
                           B(12) => A4(12), B(11) => A4(11), B(10) => A4(10), 
                           B(9) => A4(9), B(8) => A4(8), B(7) => A4(7), B(6) =>
                           A4(6), B(5) => A4(5), B(4) => A4(4), B(3) => A4(3), 
                           B(2) => A4(2), B(1) => A4(1), B(0) => A4(0), S => 
                           S(0), Y(15) => out2_15_port, Y(14) => out2_14_port, 
                           Y(13) => out2_13_port, Y(12) => out2_12_port, Y(11) 
                           => out2_11_port, Y(10) => out2_10_port, Y(9) => 
                           out2_9_port, Y(8) => out2_8_port, Y(7) => 
                           out2_7_port, Y(6) => out2_6_port, Y(5) => 
                           out2_5_port, Y(4) => out2_4_port, Y(3) => 
                           out2_3_port, Y(2) => out2_2_port, Y(1) => 
                           out2_1_port, Y(0) => out2_0_port);
   MUX3 : muxN1_N16_19 port map( A(15) => A5(15), A(14) => A5(14), A(13) => 
                           A5(13), A(12) => A5(12), A(11) => A5(11), A(10) => 
                           A5(10), A(9) => A5(9), A(8) => A5(8), A(7) => A5(7),
                           A(6) => A5(6), A(5) => A5(5), A(4) => A5(4), A(3) =>
                           A5(3), A(2) => A5(2), A(1) => A5(1), A(0) => A5(0), 
                           B(15) => A6(15), B(14) => A6(14), B(13) => A6(13), 
                           B(12) => A6(12), B(11) => A6(11), B(10) => A6(10), 
                           B(9) => A6(9), B(8) => A6(8), B(7) => A6(7), B(6) =>
                           A6(6), B(5) => A6(5), B(4) => A6(4), B(3) => A6(3), 
                           B(2) => A6(2), B(1) => A6(1), B(0) => A6(0), S => 
                           S(0), Y(15) => out3_15_port, Y(14) => out3_14_port, 
                           Y(13) => out3_13_port, Y(12) => out3_12_port, Y(11) 
                           => out3_11_port, Y(10) => out3_10_port, Y(9) => 
                           out3_9_port, Y(8) => out3_8_port, Y(7) => 
                           out3_7_port, Y(6) => out3_6_port, Y(5) => 
                           out3_5_port, Y(4) => out3_4_port, Y(3) => 
                           out3_3_port, Y(2) => out3_2_port, Y(1) => 
                           out3_1_port, Y(0) => out3_0_port);
   MUX4 : muxN1_N16_18 port map( A(15) => A7(15), A(14) => A7(14), A(13) => 
                           A7(13), A(12) => A7(12), A(11) => A7(11), A(10) => 
                           A7(10), A(9) => A7(9), A(8) => A7(8), A(7) => A7(7),
                           A(6) => A7(6), A(5) => A7(5), A(4) => A7(4), A(3) =>
                           A7(3), A(2) => A7(2), A(1) => A7(1), A(0) => A7(0), 
                           B(15) => A8(15), B(14) => A8(14), B(13) => A8(13), 
                           B(12) => A8(12), B(11) => A8(11), B(10) => A8(10), 
                           B(9) => A8(9), B(8) => A8(8), B(7) => A8(7), B(6) =>
                           A8(6), B(5) => A8(5), B(4) => A8(4), B(3) => A8(3), 
                           B(2) => A8(2), B(1) => A8(1), B(0) => A8(0), S => 
                           S(0), Y(15) => out4_15_port, Y(14) => out4_14_port, 
                           Y(13) => out4_13_port, Y(12) => out4_12_port, Y(11) 
                           => out4_11_port, Y(10) => out4_10_port, Y(9) => 
                           out4_9_port, Y(8) => out4_8_port, Y(7) => 
                           out4_7_port, Y(6) => out4_6_port, Y(5) => 
                           out4_5_port, Y(4) => out4_4_port, Y(3) => 
                           out4_3_port, Y(2) => out4_2_port, Y(1) => 
                           out4_1_port, Y(0) => out4_0_port);
   MUX5 : muxN1_N16_17 port map( A(15) => out1_15_port, A(14) => out1_14_port, 
                           A(13) => out1_13_port, A(12) => out1_12_port, A(11) 
                           => out1_11_port, A(10) => out1_10_port, A(9) => 
                           out1_9_port, A(8) => out1_8_port, A(7) => 
                           out1_7_port, A(6) => out1_6_port, A(5) => 
                           out1_5_port, A(4) => out1_4_port, A(3) => 
                           out1_3_port, A(2) => out1_2_port, A(1) => 
                           out1_1_port, A(0) => out1_0_port, B(15) => 
                           out2_15_port, B(14) => out2_14_port, B(13) => 
                           out2_13_port, B(12) => out2_12_port, B(11) => 
                           out2_11_port, B(10) => out2_10_port, B(9) => 
                           out2_9_port, B(8) => out2_8_port, B(7) => 
                           out2_7_port, B(6) => out2_6_port, B(5) => 
                           out2_5_port, B(4) => out2_4_port, B(3) => 
                           out2_3_port, B(2) => out2_2_port, B(1) => 
                           out2_1_port, B(0) => out2_0_port, S => S(1), Y(15) 
                           => out5_15_port, Y(14) => out5_14_port, Y(13) => 
                           out5_13_port, Y(12) => out5_12_port, Y(11) => 
                           out5_11_port, Y(10) => out5_10_port, Y(9) => 
                           out5_9_port, Y(8) => out5_8_port, Y(7) => 
                           out5_7_port, Y(6) => out5_6_port, Y(5) => 
                           out5_5_port, Y(4) => out5_4_port, Y(3) => 
                           out5_3_port, Y(2) => out5_2_port, Y(1) => 
                           out5_1_port, Y(0) => out5_0_port);
   MUX6 : muxN1_N16_16 port map( A(15) => out3_15_port, A(14) => out3_14_port, 
                           A(13) => out3_13_port, A(12) => out3_12_port, A(11) 
                           => out3_11_port, A(10) => out3_10_port, A(9) => 
                           out3_9_port, A(8) => out3_8_port, A(7) => 
                           out3_7_port, A(6) => out3_6_port, A(5) => 
                           out3_5_port, A(4) => out3_4_port, A(3) => 
                           out3_3_port, A(2) => out3_2_port, A(1) => 
                           out3_1_port, A(0) => out3_0_port, B(15) => 
                           out4_15_port, B(14) => out4_14_port, B(13) => 
                           out4_13_port, B(12) => out4_12_port, B(11) => 
                           out4_11_port, B(10) => out4_10_port, B(9) => 
                           out4_9_port, B(8) => out4_8_port, B(7) => 
                           out4_7_port, B(6) => out4_6_port, B(5) => 
                           out4_5_port, B(4) => out4_4_port, B(3) => 
                           out4_3_port, B(2) => out4_2_port, B(1) => 
                           out4_1_port, B(0) => out4_0_port, S => S(1), Y(15) 
                           => out6_15_port, Y(14) => out6_14_port, Y(13) => 
                           out6_13_port, Y(12) => out6_12_port, Y(11) => 
                           out6_11_port, Y(10) => out6_10_port, Y(9) => 
                           out6_9_port, Y(8) => out6_8_port, Y(7) => 
                           out6_7_port, Y(6) => out6_6_port, Y(5) => 
                           out6_5_port, Y(4) => out6_4_port, Y(3) => 
                           out6_3_port, Y(2) => out6_2_port, Y(1) => 
                           out6_1_port, Y(0) => out6_0_port);
   MUX7 : muxN1_N16_15 port map( A(15) => out5_15_port, A(14) => out5_14_port, 
                           A(13) => out5_13_port, A(12) => out5_12_port, A(11) 
                           => out5_11_port, A(10) => out5_10_port, A(9) => 
                           out5_9_port, A(8) => out5_8_port, A(7) => 
                           out5_7_port, A(6) => out5_6_port, A(5) => 
                           out5_5_port, A(4) => out5_4_port, A(3) => 
                           out5_3_port, A(2) => out5_2_port, A(1) => 
                           out5_1_port, A(0) => out5_0_port, B(15) => 
                           out6_15_port, B(14) => out6_14_port, B(13) => 
                           out6_13_port, B(12) => out6_12_port, B(11) => 
                           out6_11_port, B(10) => out6_10_port, B(9) => 
                           out6_9_port, B(8) => out6_8_port, B(7) => 
                           out6_7_port, B(6) => out6_6_port, B(5) => 
                           out6_5_port, B(4) => out6_4_port, B(3) => 
                           out6_3_port, B(2) => out6_2_port, B(1) => 
                           out6_1_port, B(0) => out6_0_port, S => S(2), Y(15) 
                           => Y(15), Y(14) => Y(14), Y(13) => Y(13), Y(12) => 
                           Y(12), Y(11) => Y(11), Y(10) => Y(10), Y(9) => Y(9),
                           Y(8) => Y(8), Y(7) => Y(7), Y(6) => Y(6), Y(5) => 
                           Y(5), Y(4) => Y(4), Y(3) => Y(3), Y(2) => Y(2), Y(1)
                           => Y(1), Y(0) => Y(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux_8to1_N16_2 is

   port( A1, A2, A3, A4, A5, A6, A7, A8 : in std_logic_vector (15 downto 0);  S
         : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end mux_8to1_N16_2;

architecture SYN_ARCHSTRUCT of mux_8to1_N16_2 is

   component muxN1_N16_8
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_9
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_10
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_11
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_12
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_13
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_14
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   signal out1_15_port, out1_14_port, out1_13_port, out1_12_port, out1_11_port,
      out1_10_port, out1_9_port, out1_8_port, out1_7_port, out1_6_port, 
      out1_5_port, out1_4_port, out1_3_port, out1_2_port, out1_1_port, 
      out1_0_port, out2_15_port, out2_14_port, out2_13_port, out2_12_port, 
      out2_11_port, out2_10_port, out2_9_port, out2_8_port, out2_7_port, 
      out2_6_port, out2_5_port, out2_4_port, out2_3_port, out2_2_port, 
      out2_1_port, out2_0_port, out3_15_port, out3_14_port, out3_13_port, 
      out3_12_port, out3_11_port, out3_10_port, out3_9_port, out3_8_port, 
      out3_7_port, out3_6_port, out3_5_port, out3_4_port, out3_3_port, 
      out3_2_port, out3_1_port, out3_0_port, out4_15_port, out4_14_port, 
      out4_13_port, out4_12_port, out4_11_port, out4_10_port, out4_9_port, 
      out4_8_port, out4_7_port, out4_6_port, out4_5_port, out4_4_port, 
      out4_3_port, out4_2_port, out4_1_port, out4_0_port, out5_15_port, 
      out5_14_port, out5_13_port, out5_12_port, out5_11_port, out5_10_port, 
      out5_9_port, out5_8_port, out5_7_port, out5_6_port, out5_5_port, 
      out5_4_port, out5_3_port, out5_2_port, out5_1_port, out5_0_port, 
      out6_15_port, out6_14_port, out6_13_port, out6_12_port, out6_11_port, 
      out6_10_port, out6_9_port, out6_8_port, out6_7_port, out6_6_port, 
      out6_5_port, out6_4_port, out6_3_port, out6_2_port, out6_1_port, 
      out6_0_port : std_logic;

begin
   
   MUX1 : muxN1_N16_14 port map( A(15) => A1(15), A(14) => A1(14), A(13) => 
                           A1(13), A(12) => A1(12), A(11) => A1(11), A(10) => 
                           A1(10), A(9) => A1(9), A(8) => A1(8), A(7) => A1(7),
                           A(6) => A1(6), A(5) => A1(5), A(4) => A1(4), A(3) =>
                           A1(3), A(2) => A1(2), A(1) => A1(1), A(0) => A1(0), 
                           B(15) => A2(15), B(14) => A2(14), B(13) => A2(13), 
                           B(12) => A2(12), B(11) => A2(11), B(10) => A2(10), 
                           B(9) => A2(9), B(8) => A2(8), B(7) => A2(7), B(6) =>
                           A2(6), B(5) => A2(5), B(4) => A2(4), B(3) => A2(3), 
                           B(2) => A2(2), B(1) => A2(1), B(0) => A2(0), S => 
                           S(0), Y(15) => out1_15_port, Y(14) => out1_14_port, 
                           Y(13) => out1_13_port, Y(12) => out1_12_port, Y(11) 
                           => out1_11_port, Y(10) => out1_10_port, Y(9) => 
                           out1_9_port, Y(8) => out1_8_port, Y(7) => 
                           out1_7_port, Y(6) => out1_6_port, Y(5) => 
                           out1_5_port, Y(4) => out1_4_port, Y(3) => 
                           out1_3_port, Y(2) => out1_2_port, Y(1) => 
                           out1_1_port, Y(0) => out1_0_port);
   MUX2 : muxN1_N16_13 port map( A(15) => A3(15), A(14) => A3(14), A(13) => 
                           A3(13), A(12) => A3(12), A(11) => A3(11), A(10) => 
                           A3(10), A(9) => A3(9), A(8) => A3(8), A(7) => A3(7),
                           A(6) => A3(6), A(5) => A3(5), A(4) => A3(4), A(3) =>
                           A3(3), A(2) => A3(2), A(1) => A3(1), A(0) => A3(0), 
                           B(15) => A4(15), B(14) => A4(14), B(13) => A4(13), 
                           B(12) => A4(12), B(11) => A4(11), B(10) => A4(10), 
                           B(9) => A4(9), B(8) => A4(8), B(7) => A4(7), B(6) =>
                           A4(6), B(5) => A4(5), B(4) => A4(4), B(3) => A4(3), 
                           B(2) => A4(2), B(1) => A4(1), B(0) => A4(0), S => 
                           S(0), Y(15) => out2_15_port, Y(14) => out2_14_port, 
                           Y(13) => out2_13_port, Y(12) => out2_12_port, Y(11) 
                           => out2_11_port, Y(10) => out2_10_port, Y(9) => 
                           out2_9_port, Y(8) => out2_8_port, Y(7) => 
                           out2_7_port, Y(6) => out2_6_port, Y(5) => 
                           out2_5_port, Y(4) => out2_4_port, Y(3) => 
                           out2_3_port, Y(2) => out2_2_port, Y(1) => 
                           out2_1_port, Y(0) => out2_0_port);
   MUX3 : muxN1_N16_12 port map( A(15) => A5(15), A(14) => A5(14), A(13) => 
                           A5(13), A(12) => A5(12), A(11) => A5(11), A(10) => 
                           A5(10), A(9) => A5(9), A(8) => A5(8), A(7) => A5(7),
                           A(6) => A5(6), A(5) => A5(5), A(4) => A5(4), A(3) =>
                           A5(3), A(2) => A5(2), A(1) => A5(1), A(0) => A5(0), 
                           B(15) => A6(15), B(14) => A6(14), B(13) => A6(13), 
                           B(12) => A6(12), B(11) => A6(11), B(10) => A6(10), 
                           B(9) => A6(9), B(8) => A6(8), B(7) => A6(7), B(6) =>
                           A6(6), B(5) => A6(5), B(4) => A6(4), B(3) => A6(3), 
                           B(2) => A6(2), B(1) => A6(1), B(0) => A6(0), S => 
                           S(0), Y(15) => out3_15_port, Y(14) => out3_14_port, 
                           Y(13) => out3_13_port, Y(12) => out3_12_port, Y(11) 
                           => out3_11_port, Y(10) => out3_10_port, Y(9) => 
                           out3_9_port, Y(8) => out3_8_port, Y(7) => 
                           out3_7_port, Y(6) => out3_6_port, Y(5) => 
                           out3_5_port, Y(4) => out3_4_port, Y(3) => 
                           out3_3_port, Y(2) => out3_2_port, Y(1) => 
                           out3_1_port, Y(0) => out3_0_port);
   MUX4 : muxN1_N16_11 port map( A(15) => A7(15), A(14) => A7(14), A(13) => 
                           A7(13), A(12) => A7(12), A(11) => A7(11), A(10) => 
                           A7(10), A(9) => A7(9), A(8) => A7(8), A(7) => A7(7),
                           A(6) => A7(6), A(5) => A7(5), A(4) => A7(4), A(3) =>
                           A7(3), A(2) => A7(2), A(1) => A7(1), A(0) => A7(0), 
                           B(15) => A8(15), B(14) => A8(14), B(13) => A8(13), 
                           B(12) => A8(12), B(11) => A8(11), B(10) => A8(10), 
                           B(9) => A8(9), B(8) => A8(8), B(7) => A8(7), B(6) =>
                           A8(6), B(5) => A8(5), B(4) => A8(4), B(3) => A8(3), 
                           B(2) => A8(2), B(1) => A8(1), B(0) => A8(0), S => 
                           S(0), Y(15) => out4_15_port, Y(14) => out4_14_port, 
                           Y(13) => out4_13_port, Y(12) => out4_12_port, Y(11) 
                           => out4_11_port, Y(10) => out4_10_port, Y(9) => 
                           out4_9_port, Y(8) => out4_8_port, Y(7) => 
                           out4_7_port, Y(6) => out4_6_port, Y(5) => 
                           out4_5_port, Y(4) => out4_4_port, Y(3) => 
                           out4_3_port, Y(2) => out4_2_port, Y(1) => 
                           out4_1_port, Y(0) => out4_0_port);
   MUX5 : muxN1_N16_10 port map( A(15) => out1_15_port, A(14) => out1_14_port, 
                           A(13) => out1_13_port, A(12) => out1_12_port, A(11) 
                           => out1_11_port, A(10) => out1_10_port, A(9) => 
                           out1_9_port, A(8) => out1_8_port, A(7) => 
                           out1_7_port, A(6) => out1_6_port, A(5) => 
                           out1_5_port, A(4) => out1_4_port, A(3) => 
                           out1_3_port, A(2) => out1_2_port, A(1) => 
                           out1_1_port, A(0) => out1_0_port, B(15) => 
                           out2_15_port, B(14) => out2_14_port, B(13) => 
                           out2_13_port, B(12) => out2_12_port, B(11) => 
                           out2_11_port, B(10) => out2_10_port, B(9) => 
                           out2_9_port, B(8) => out2_8_port, B(7) => 
                           out2_7_port, B(6) => out2_6_port, B(5) => 
                           out2_5_port, B(4) => out2_4_port, B(3) => 
                           out2_3_port, B(2) => out2_2_port, B(1) => 
                           out2_1_port, B(0) => out2_0_port, S => S(1), Y(15) 
                           => out5_15_port, Y(14) => out5_14_port, Y(13) => 
                           out5_13_port, Y(12) => out5_12_port, Y(11) => 
                           out5_11_port, Y(10) => out5_10_port, Y(9) => 
                           out5_9_port, Y(8) => out5_8_port, Y(7) => 
                           out5_7_port, Y(6) => out5_6_port, Y(5) => 
                           out5_5_port, Y(4) => out5_4_port, Y(3) => 
                           out5_3_port, Y(2) => out5_2_port, Y(1) => 
                           out5_1_port, Y(0) => out5_0_port);
   MUX6 : muxN1_N16_9 port map( A(15) => out3_15_port, A(14) => out3_14_port, 
                           A(13) => out3_13_port, A(12) => out3_12_port, A(11) 
                           => out3_11_port, A(10) => out3_10_port, A(9) => 
                           out3_9_port, A(8) => out3_8_port, A(7) => 
                           out3_7_port, A(6) => out3_6_port, A(5) => 
                           out3_5_port, A(4) => out3_4_port, A(3) => 
                           out3_3_port, A(2) => out3_2_port, A(1) => 
                           out3_1_port, A(0) => out3_0_port, B(15) => 
                           out4_15_port, B(14) => out4_14_port, B(13) => 
                           out4_13_port, B(12) => out4_12_port, B(11) => 
                           out4_11_port, B(10) => out4_10_port, B(9) => 
                           out4_9_port, B(8) => out4_8_port, B(7) => 
                           out4_7_port, B(6) => out4_6_port, B(5) => 
                           out4_5_port, B(4) => out4_4_port, B(3) => 
                           out4_3_port, B(2) => out4_2_port, B(1) => 
                           out4_1_port, B(0) => out4_0_port, S => S(1), Y(15) 
                           => out6_15_port, Y(14) => out6_14_port, Y(13) => 
                           out6_13_port, Y(12) => out6_12_port, Y(11) => 
                           out6_11_port, Y(10) => out6_10_port, Y(9) => 
                           out6_9_port, Y(8) => out6_8_port, Y(7) => 
                           out6_7_port, Y(6) => out6_6_port, Y(5) => 
                           out6_5_port, Y(4) => out6_4_port, Y(3) => 
                           out6_3_port, Y(2) => out6_2_port, Y(1) => 
                           out6_1_port, Y(0) => out6_0_port);
   MUX7 : muxN1_N16_8 port map( A(15) => out5_15_port, A(14) => out5_14_port, 
                           A(13) => out5_13_port, A(12) => out5_12_port, A(11) 
                           => out5_11_port, A(10) => out5_10_port, A(9) => 
                           out5_9_port, A(8) => out5_8_port, A(7) => 
                           out5_7_port, A(6) => out5_6_port, A(5) => 
                           out5_5_port, A(4) => out5_4_port, A(3) => 
                           out5_3_port, A(2) => out5_2_port, A(1) => 
                           out5_1_port, A(0) => out5_0_port, B(15) => 
                           out6_15_port, B(14) => out6_14_port, B(13) => 
                           out6_13_port, B(12) => out6_12_port, B(11) => 
                           out6_11_port, B(10) => out6_10_port, B(9) => 
                           out6_9_port, B(8) => out6_8_port, B(7) => 
                           out6_7_port, B(6) => out6_6_port, B(5) => 
                           out6_5_port, B(4) => out6_4_port, B(3) => 
                           out6_3_port, B(2) => out6_2_port, B(1) => 
                           out6_1_port, B(0) => out6_0_port, S => S(2), Y(15) 
                           => Y(15), Y(14) => Y(14), Y(13) => Y(13), Y(12) => 
                           Y(12), Y(11) => Y(11), Y(10) => Y(10), Y(9) => Y(9),
                           Y(8) => Y(8), Y(7) => Y(7), Y(6) => Y(6), Y(5) => 
                           Y(5), Y(4) => Y(4), Y(3) => Y(3), Y(2) => Y(2), Y(1)
                           => Y(1), Y(0) => Y(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux_8to1_N16_1 is

   port( A1, A2, A3, A4, A5, A6, A7, A8 : in std_logic_vector (15 downto 0);  S
         : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end mux_8to1_N16_1;

architecture SYN_ARCHSTRUCT of mux_8to1_N16_1 is

   component muxN1_N16_1
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_2
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_3
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_4
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_5
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_6
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_7
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   signal out1_15_port, out1_14_port, out1_13_port, out1_12_port, out1_11_port,
      out1_10_port, out1_9_port, out1_8_port, out1_7_port, out1_6_port, 
      out1_5_port, out1_4_port, out1_3_port, out1_2_port, out1_1_port, 
      out1_0_port, out2_15_port, out2_14_port, out2_13_port, out2_12_port, 
      out2_11_port, out2_10_port, out2_9_port, out2_8_port, out2_7_port, 
      out2_6_port, out2_5_port, out2_4_port, out2_3_port, out2_2_port, 
      out2_1_port, out2_0_port, out3_15_port, out3_14_port, out3_13_port, 
      out3_12_port, out3_11_port, out3_10_port, out3_9_port, out3_8_port, 
      out3_7_port, out3_6_port, out3_5_port, out3_4_port, out3_3_port, 
      out3_2_port, out3_1_port, out3_0_port, out4_15_port, out4_14_port, 
      out4_13_port, out4_12_port, out4_11_port, out4_10_port, out4_9_port, 
      out4_8_port, out4_7_port, out4_6_port, out4_5_port, out4_4_port, 
      out4_3_port, out4_2_port, out4_1_port, out4_0_port, out5_15_port, 
      out5_14_port, out5_13_port, out5_12_port, out5_11_port, out5_10_port, 
      out5_9_port, out5_8_port, out5_7_port, out5_6_port, out5_5_port, 
      out5_4_port, out5_3_port, out5_2_port, out5_1_port, out5_0_port, 
      out6_15_port, out6_14_port, out6_13_port, out6_12_port, out6_11_port, 
      out6_10_port, out6_9_port, out6_8_port, out6_7_port, out6_6_port, 
      out6_5_port, out6_4_port, out6_3_port, out6_2_port, out6_1_port, 
      out6_0_port : std_logic;

begin
   
   MUX1 : muxN1_N16_7 port map( A(15) => A1(15), A(14) => A1(14), A(13) => 
                           A1(13), A(12) => A1(12), A(11) => A1(11), A(10) => 
                           A1(10), A(9) => A1(9), A(8) => A1(8), A(7) => A1(7),
                           A(6) => A1(6), A(5) => A1(5), A(4) => A1(4), A(3) =>
                           A1(3), A(2) => A1(2), A(1) => A1(1), A(0) => A1(0), 
                           B(15) => A2(15), B(14) => A2(14), B(13) => A2(13), 
                           B(12) => A2(12), B(11) => A2(11), B(10) => A2(10), 
                           B(9) => A2(9), B(8) => A2(8), B(7) => A2(7), B(6) =>
                           A2(6), B(5) => A2(5), B(4) => A2(4), B(3) => A2(3), 
                           B(2) => A2(2), B(1) => A2(1), B(0) => A2(0), S => 
                           S(0), Y(15) => out1_15_port, Y(14) => out1_14_port, 
                           Y(13) => out1_13_port, Y(12) => out1_12_port, Y(11) 
                           => out1_11_port, Y(10) => out1_10_port, Y(9) => 
                           out1_9_port, Y(8) => out1_8_port, Y(7) => 
                           out1_7_port, Y(6) => out1_6_port, Y(5) => 
                           out1_5_port, Y(4) => out1_4_port, Y(3) => 
                           out1_3_port, Y(2) => out1_2_port, Y(1) => 
                           out1_1_port, Y(0) => out1_0_port);
   MUX2 : muxN1_N16_6 port map( A(15) => A3(15), A(14) => A3(14), A(13) => 
                           A3(13), A(12) => A3(12), A(11) => A3(11), A(10) => 
                           A3(10), A(9) => A3(9), A(8) => A3(8), A(7) => A3(7),
                           A(6) => A3(6), A(5) => A3(5), A(4) => A3(4), A(3) =>
                           A3(3), A(2) => A3(2), A(1) => A3(1), A(0) => A3(0), 
                           B(15) => A4(15), B(14) => A4(14), B(13) => A4(13), 
                           B(12) => A4(12), B(11) => A4(11), B(10) => A4(10), 
                           B(9) => A4(9), B(8) => A4(8), B(7) => A4(7), B(6) =>
                           A4(6), B(5) => A4(5), B(4) => A4(4), B(3) => A4(3), 
                           B(2) => A4(2), B(1) => A4(1), B(0) => A4(0), S => 
                           S(0), Y(15) => out2_15_port, Y(14) => out2_14_port, 
                           Y(13) => out2_13_port, Y(12) => out2_12_port, Y(11) 
                           => out2_11_port, Y(10) => out2_10_port, Y(9) => 
                           out2_9_port, Y(8) => out2_8_port, Y(7) => 
                           out2_7_port, Y(6) => out2_6_port, Y(5) => 
                           out2_5_port, Y(4) => out2_4_port, Y(3) => 
                           out2_3_port, Y(2) => out2_2_port, Y(1) => 
                           out2_1_port, Y(0) => out2_0_port);
   MUX3 : muxN1_N16_5 port map( A(15) => A5(15), A(14) => A5(14), A(13) => 
                           A5(13), A(12) => A5(12), A(11) => A5(11), A(10) => 
                           A5(10), A(9) => A5(9), A(8) => A5(8), A(7) => A5(7),
                           A(6) => A5(6), A(5) => A5(5), A(4) => A5(4), A(3) =>
                           A5(3), A(2) => A5(2), A(1) => A5(1), A(0) => A5(0), 
                           B(15) => A6(15), B(14) => A6(14), B(13) => A6(13), 
                           B(12) => A6(12), B(11) => A6(11), B(10) => A6(10), 
                           B(9) => A6(9), B(8) => A6(8), B(7) => A6(7), B(6) =>
                           A6(6), B(5) => A6(5), B(4) => A6(4), B(3) => A6(3), 
                           B(2) => A6(2), B(1) => A6(1), B(0) => A6(0), S => 
                           S(0), Y(15) => out3_15_port, Y(14) => out3_14_port, 
                           Y(13) => out3_13_port, Y(12) => out3_12_port, Y(11) 
                           => out3_11_port, Y(10) => out3_10_port, Y(9) => 
                           out3_9_port, Y(8) => out3_8_port, Y(7) => 
                           out3_7_port, Y(6) => out3_6_port, Y(5) => 
                           out3_5_port, Y(4) => out3_4_port, Y(3) => 
                           out3_3_port, Y(2) => out3_2_port, Y(1) => 
                           out3_1_port, Y(0) => out3_0_port);
   MUX4 : muxN1_N16_4 port map( A(15) => A7(15), A(14) => A7(14), A(13) => 
                           A7(13), A(12) => A7(12), A(11) => A7(11), A(10) => 
                           A7(10), A(9) => A7(9), A(8) => A7(8), A(7) => A7(7),
                           A(6) => A7(6), A(5) => A7(5), A(4) => A7(4), A(3) =>
                           A7(3), A(2) => A7(2), A(1) => A7(1), A(0) => A7(0), 
                           B(15) => A8(15), B(14) => A8(14), B(13) => A8(13), 
                           B(12) => A8(12), B(11) => A8(11), B(10) => A8(10), 
                           B(9) => A8(9), B(8) => A8(8), B(7) => A8(7), B(6) =>
                           A8(6), B(5) => A8(5), B(4) => A8(4), B(3) => A8(3), 
                           B(2) => A8(2), B(1) => A8(1), B(0) => A8(0), S => 
                           S(0), Y(15) => out4_15_port, Y(14) => out4_14_port, 
                           Y(13) => out4_13_port, Y(12) => out4_12_port, Y(11) 
                           => out4_11_port, Y(10) => out4_10_port, Y(9) => 
                           out4_9_port, Y(8) => out4_8_port, Y(7) => 
                           out4_7_port, Y(6) => out4_6_port, Y(5) => 
                           out4_5_port, Y(4) => out4_4_port, Y(3) => 
                           out4_3_port, Y(2) => out4_2_port, Y(1) => 
                           out4_1_port, Y(0) => out4_0_port);
   MUX5 : muxN1_N16_3 port map( A(15) => out1_15_port, A(14) => out1_14_port, 
                           A(13) => out1_13_port, A(12) => out1_12_port, A(11) 
                           => out1_11_port, A(10) => out1_10_port, A(9) => 
                           out1_9_port, A(8) => out1_8_port, A(7) => 
                           out1_7_port, A(6) => out1_6_port, A(5) => 
                           out1_5_port, A(4) => out1_4_port, A(3) => 
                           out1_3_port, A(2) => out1_2_port, A(1) => 
                           out1_1_port, A(0) => out1_0_port, B(15) => 
                           out2_15_port, B(14) => out2_14_port, B(13) => 
                           out2_13_port, B(12) => out2_12_port, B(11) => 
                           out2_11_port, B(10) => out2_10_port, B(9) => 
                           out2_9_port, B(8) => out2_8_port, B(7) => 
                           out2_7_port, B(6) => out2_6_port, B(5) => 
                           out2_5_port, B(4) => out2_4_port, B(3) => 
                           out2_3_port, B(2) => out2_2_port, B(1) => 
                           out2_1_port, B(0) => out2_0_port, S => S(1), Y(15) 
                           => out5_15_port, Y(14) => out5_14_port, Y(13) => 
                           out5_13_port, Y(12) => out5_12_port, Y(11) => 
                           out5_11_port, Y(10) => out5_10_port, Y(9) => 
                           out5_9_port, Y(8) => out5_8_port, Y(7) => 
                           out5_7_port, Y(6) => out5_6_port, Y(5) => 
                           out5_5_port, Y(4) => out5_4_port, Y(3) => 
                           out5_3_port, Y(2) => out5_2_port, Y(1) => 
                           out5_1_port, Y(0) => out5_0_port);
   MUX6 : muxN1_N16_2 port map( A(15) => out3_15_port, A(14) => out3_14_port, 
                           A(13) => out3_13_port, A(12) => out3_12_port, A(11) 
                           => out3_11_port, A(10) => out3_10_port, A(9) => 
                           out3_9_port, A(8) => out3_8_port, A(7) => 
                           out3_7_port, A(6) => out3_6_port, A(5) => 
                           out3_5_port, A(4) => out3_4_port, A(3) => 
                           out3_3_port, A(2) => out3_2_port, A(1) => 
                           out3_1_port, A(0) => out3_0_port, B(15) => 
                           out4_15_port, B(14) => out4_14_port, B(13) => 
                           out4_13_port, B(12) => out4_12_port, B(11) => 
                           out4_11_port, B(10) => out4_10_port, B(9) => 
                           out4_9_port, B(8) => out4_8_port, B(7) => 
                           out4_7_port, B(6) => out4_6_port, B(5) => 
                           out4_5_port, B(4) => out4_4_port, B(3) => 
                           out4_3_port, B(2) => out4_2_port, B(1) => 
                           out4_1_port, B(0) => out4_0_port, S => S(1), Y(15) 
                           => out6_15_port, Y(14) => out6_14_port, Y(13) => 
                           out6_13_port, Y(12) => out6_12_port, Y(11) => 
                           out6_11_port, Y(10) => out6_10_port, Y(9) => 
                           out6_9_port, Y(8) => out6_8_port, Y(7) => 
                           out6_7_port, Y(6) => out6_6_port, Y(5) => 
                           out6_5_port, Y(4) => out6_4_port, Y(3) => 
                           out6_3_port, Y(2) => out6_2_port, Y(1) => 
                           out6_1_port, Y(0) => out6_0_port);
   MUX7 : muxN1_N16_1 port map( A(15) => out5_15_port, A(14) => out5_14_port, 
                           A(13) => out5_13_port, A(12) => out5_12_port, A(11) 
                           => out5_11_port, A(10) => out5_10_port, A(9) => 
                           out5_9_port, A(8) => out5_8_port, A(7) => 
                           out5_7_port, A(6) => out5_6_port, A(5) => 
                           out5_5_port, A(4) => out5_4_port, A(3) => 
                           out5_3_port, A(2) => out5_2_port, A(1) => 
                           out5_1_port, A(0) => out5_0_port, B(15) => 
                           out6_15_port, B(14) => out6_14_port, B(13) => 
                           out6_13_port, B(12) => out6_12_port, B(11) => 
                           out6_11_port, B(10) => out6_10_port, B(9) => 
                           out6_9_port, B(8) => out6_8_port, B(7) => 
                           out6_7_port, B(6) => out6_6_port, B(5) => 
                           out6_5_port, B(4) => out6_4_port, B(3) => 
                           out6_3_port, B(2) => out6_2_port, B(1) => 
                           out6_1_port, B(0) => out6_0_port, S => S(2), Y(15) 
                           => Y(15), Y(14) => Y(14), Y(13) => Y(13), Y(12) => 
                           Y(12), Y(11) => Y(11), Y(10) => Y(10), Y(9) => Y(9),
                           Y(8) => Y(8), Y(7) => Y(7), Y(6) => Y(6), Y(5) => 
                           Y(5), Y(4) => Y(4), Y(3) => Y(3), Y(2) => Y(2), Y(1)
                           => Y(1), Y(0) => Y(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_7 is

   port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end complementor_N16_7;

architecture SYN_ARCHDATAFLOW of complementor_N16_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component complementor_N16_7_DW01_inc_0_DW01_inc_6
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal N9, N8, N7, N6, N5, N4, N3, N2, N15, N14, N13, N12, N11, N10, N1, N0 
      : std_logic;

begin
   
   add_0_root_add_19_ni : complementor_N16_7_DW01_inc_0_DW01_inc_6 port map( 
                           A(15) => N0, A(14) => N1, A(13) => N2, A(12) => N3, 
                           A(11) => N4, A(10) => N5, A(9) => N6, A(8) => N7, 
                           A(7) => N8, A(6) => N9, A(5) => N10, A(4) => N11, 
                           A(3) => N12, A(2) => N13, A(1) => N14, A(0) => N15, 
                           SUM(15) => Y(15), SUM(14) => Y(14), SUM(13) => Y(13)
                           , SUM(12) => Y(12), SUM(11) => Y(11), SUM(10) => 
                           Y(10), SUM(9) => Y(9), SUM(8) => Y(8), SUM(7) => 
                           Y(7), SUM(6) => Y(6), SUM(5) => Y(5), SUM(4) => Y(4)
                           , SUM(3) => Y(3), SUM(2) => Y(2), SUM(1) => Y(1), 
                           SUM(0) => Y(0));
   U2 : INV_X1 port map( A => A(6), ZN => N9);
   U3 : INV_X1 port map( A => A(7), ZN => N8);
   U4 : INV_X1 port map( A => A(8), ZN => N7);
   U5 : INV_X1 port map( A => A(9), ZN => N6);
   U6 : INV_X1 port map( A => A(10), ZN => N5);
   U7 : INV_X1 port map( A => A(11), ZN => N4);
   U8 : INV_X1 port map( A => A(12), ZN => N3);
   U9 : INV_X1 port map( A => A(13), ZN => N2);
   U10 : INV_X1 port map( A => A(0), ZN => N15);
   U11 : INV_X1 port map( A => A(1), ZN => N14);
   U12 : INV_X1 port map( A => A(2), ZN => N13);
   U13 : INV_X1 port map( A => A(3), ZN => N12);
   U14 : INV_X1 port map( A => A(4), ZN => N11);
   U15 : INV_X1 port map( A => A(5), ZN => N10);
   U16 : INV_X1 port map( A => A(14), ZN => N1);
   U17 : INV_X1 port map( A => A(15), ZN => N0);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_6 is

   port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end complementor_N16_6;

architecture SYN_ARCHDATAFLOW of complementor_N16_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component complementor_N16_6_DW01_inc_0_DW01_inc_5
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal N9, N8, N7, N6, N5, N4, N3, N2, N15, N14, N13, N12, N11, N10, N1, N0 
      : std_logic;

begin
   
   add_0_root_add_19_ni : complementor_N16_6_DW01_inc_0_DW01_inc_5 port map( 
                           A(15) => N0, A(14) => N1, A(13) => N2, A(12) => N3, 
                           A(11) => N4, A(10) => N5, A(9) => N6, A(8) => N7, 
                           A(7) => N8, A(6) => N9, A(5) => N10, A(4) => N11, 
                           A(3) => N12, A(2) => N13, A(1) => N14, A(0) => N15, 
                           SUM(15) => Y(15), SUM(14) => Y(14), SUM(13) => Y(13)
                           , SUM(12) => Y(12), SUM(11) => Y(11), SUM(10) => 
                           Y(10), SUM(9) => Y(9), SUM(8) => Y(8), SUM(7) => 
                           Y(7), SUM(6) => Y(6), SUM(5) => Y(5), SUM(4) => Y(4)
                           , SUM(3) => Y(3), SUM(2) => Y(2), SUM(1) => Y(1), 
                           SUM(0) => Y(0));
   U2 : INV_X1 port map( A => A(6), ZN => N9);
   U3 : INV_X1 port map( A => A(7), ZN => N8);
   U4 : INV_X1 port map( A => A(8), ZN => N7);
   U5 : INV_X1 port map( A => A(9), ZN => N6);
   U6 : INV_X1 port map( A => A(10), ZN => N5);
   U7 : INV_X1 port map( A => A(11), ZN => N4);
   U8 : INV_X1 port map( A => A(12), ZN => N3);
   U9 : INV_X1 port map( A => A(13), ZN => N2);
   U10 : INV_X1 port map( A => A(0), ZN => N15);
   U11 : INV_X1 port map( A => A(1), ZN => N14);
   U12 : INV_X1 port map( A => A(2), ZN => N13);
   U13 : INV_X1 port map( A => A(3), ZN => N12);
   U14 : INV_X1 port map( A => A(4), ZN => N11);
   U15 : INV_X1 port map( A => A(5), ZN => N10);
   U16 : INV_X1 port map( A => A(14), ZN => N1);
   U17 : INV_X1 port map( A => A(15), ZN => N0);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_5 is

   port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end complementor_N16_5;

architecture SYN_ARCHDATAFLOW of complementor_N16_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component complementor_N16_5_DW01_inc_0_DW01_inc_4
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal N9, N8, N7, N6, N5, N4, N3, N2, N15, N14, N13, N12, N11, N10, N1, N0 
      : std_logic;

begin
   
   add_0_root_add_19_ni : complementor_N16_5_DW01_inc_0_DW01_inc_4 port map( 
                           A(15) => N0, A(14) => N1, A(13) => N2, A(12) => N3, 
                           A(11) => N4, A(10) => N5, A(9) => N6, A(8) => N7, 
                           A(7) => N8, A(6) => N9, A(5) => N10, A(4) => N11, 
                           A(3) => N12, A(2) => N13, A(1) => N14, A(0) => N15, 
                           SUM(15) => Y(15), SUM(14) => Y(14), SUM(13) => Y(13)
                           , SUM(12) => Y(12), SUM(11) => Y(11), SUM(10) => 
                           Y(10), SUM(9) => Y(9), SUM(8) => Y(8), SUM(7) => 
                           Y(7), SUM(6) => Y(6), SUM(5) => Y(5), SUM(4) => Y(4)
                           , SUM(3) => Y(3), SUM(2) => Y(2), SUM(1) => Y(1), 
                           SUM(0) => Y(0));
   U2 : INV_X1 port map( A => A(6), ZN => N9);
   U3 : INV_X1 port map( A => A(7), ZN => N8);
   U4 : INV_X1 port map( A => A(8), ZN => N7);
   U5 : INV_X1 port map( A => A(9), ZN => N6);
   U6 : INV_X1 port map( A => A(10), ZN => N5);
   U7 : INV_X1 port map( A => A(11), ZN => N4);
   U8 : INV_X1 port map( A => A(12), ZN => N3);
   U9 : INV_X1 port map( A => A(13), ZN => N2);
   U10 : INV_X1 port map( A => A(0), ZN => N15);
   U11 : INV_X1 port map( A => A(1), ZN => N14);
   U12 : INV_X1 port map( A => A(2), ZN => N13);
   U13 : INV_X1 port map( A => A(3), ZN => N12);
   U14 : INV_X1 port map( A => A(4), ZN => N11);
   U15 : INV_X1 port map( A => A(5), ZN => N10);
   U16 : INV_X1 port map( A => A(14), ZN => N1);
   U17 : INV_X1 port map( A => A(15), ZN => N0);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_4 is

   port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end complementor_N16_4;

architecture SYN_ARCHDATAFLOW of complementor_N16_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component complementor_N16_4_DW01_inc_0_DW01_inc_3
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal N9, N8, N7, N6, N5, N4, N3, N2, N15, N14, N13, N12, N11, N10, N1, N0 
      : std_logic;

begin
   
   add_0_root_add_19_ni : complementor_N16_4_DW01_inc_0_DW01_inc_3 port map( 
                           A(15) => N0, A(14) => N1, A(13) => N2, A(12) => N3, 
                           A(11) => N4, A(10) => N5, A(9) => N6, A(8) => N7, 
                           A(7) => N8, A(6) => N9, A(5) => N10, A(4) => N11, 
                           A(3) => N12, A(2) => N13, A(1) => N14, A(0) => N15, 
                           SUM(15) => Y(15), SUM(14) => Y(14), SUM(13) => Y(13)
                           , SUM(12) => Y(12), SUM(11) => Y(11), SUM(10) => 
                           Y(10), SUM(9) => Y(9), SUM(8) => Y(8), SUM(7) => 
                           Y(7), SUM(6) => Y(6), SUM(5) => Y(5), SUM(4) => Y(4)
                           , SUM(3) => Y(3), SUM(2) => Y(2), SUM(1) => Y(1), 
                           SUM(0) => Y(0));
   U2 : INV_X1 port map( A => A(6), ZN => N9);
   U3 : INV_X1 port map( A => A(7), ZN => N8);
   U4 : INV_X1 port map( A => A(8), ZN => N7);
   U5 : INV_X1 port map( A => A(9), ZN => N6);
   U6 : INV_X1 port map( A => A(10), ZN => N5);
   U7 : INV_X1 port map( A => A(11), ZN => N4);
   U8 : INV_X1 port map( A => A(12), ZN => N3);
   U9 : INV_X1 port map( A => A(13), ZN => N2);
   U10 : INV_X1 port map( A => A(0), ZN => N15);
   U11 : INV_X1 port map( A => A(1), ZN => N14);
   U12 : INV_X1 port map( A => A(2), ZN => N13);
   U13 : INV_X1 port map( A => A(3), ZN => N12);
   U14 : INV_X1 port map( A => A(4), ZN => N11);
   U15 : INV_X1 port map( A => A(5), ZN => N10);
   U16 : INV_X1 port map( A => A(14), ZN => N1);
   U17 : INV_X1 port map( A => A(15), ZN => N0);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_3 is

   port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end complementor_N16_3;

architecture SYN_ARCHDATAFLOW of complementor_N16_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component complementor_N16_3_DW01_inc_0_DW01_inc_2
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal N9, N8, N7, N6, N5, N4, N3, N2, N15, N14, N13, N12, N11, N10, N1, N0 
      : std_logic;

begin
   
   add_0_root_add_19_ni : complementor_N16_3_DW01_inc_0_DW01_inc_2 port map( 
                           A(15) => N0, A(14) => N1, A(13) => N2, A(12) => N3, 
                           A(11) => N4, A(10) => N5, A(9) => N6, A(8) => N7, 
                           A(7) => N8, A(6) => N9, A(5) => N10, A(4) => N11, 
                           A(3) => N12, A(2) => N13, A(1) => N14, A(0) => N15, 
                           SUM(15) => Y(15), SUM(14) => Y(14), SUM(13) => Y(13)
                           , SUM(12) => Y(12), SUM(11) => Y(11), SUM(10) => 
                           Y(10), SUM(9) => Y(9), SUM(8) => Y(8), SUM(7) => 
                           Y(7), SUM(6) => Y(6), SUM(5) => Y(5), SUM(4) => Y(4)
                           , SUM(3) => Y(3), SUM(2) => Y(2), SUM(1) => Y(1), 
                           SUM(0) => Y(0));
   U2 : INV_X1 port map( A => A(6), ZN => N9);
   U3 : INV_X1 port map( A => A(7), ZN => N8);
   U4 : INV_X1 port map( A => A(8), ZN => N7);
   U5 : INV_X1 port map( A => A(9), ZN => N6);
   U6 : INV_X1 port map( A => A(10), ZN => N5);
   U7 : INV_X1 port map( A => A(11), ZN => N4);
   U8 : INV_X1 port map( A => A(12), ZN => N3);
   U9 : INV_X1 port map( A => A(13), ZN => N2);
   U10 : INV_X1 port map( A => A(0), ZN => N15);
   U11 : INV_X1 port map( A => A(1), ZN => N14);
   U12 : INV_X1 port map( A => A(2), ZN => N13);
   U13 : INV_X1 port map( A => A(3), ZN => N12);
   U14 : INV_X1 port map( A => A(4), ZN => N11);
   U15 : INV_X1 port map( A => A(5), ZN => N10);
   U16 : INV_X1 port map( A => A(14), ZN => N1);
   U17 : INV_X1 port map( A => A(15), ZN => N0);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_2 is

   port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end complementor_N16_2;

architecture SYN_ARCHDATAFLOW of complementor_N16_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component complementor_N16_2_DW01_inc_0_DW01_inc_1
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal N9, N8, N7, N6, N5, N4, N3, N2, N15, N14, N13, N12, N11, N10, N1, N0 
      : std_logic;

begin
   
   add_0_root_add_19_ni : complementor_N16_2_DW01_inc_0_DW01_inc_1 port map( 
                           A(15) => N0, A(14) => N1, A(13) => N2, A(12) => N3, 
                           A(11) => N4, A(10) => N5, A(9) => N6, A(8) => N7, 
                           A(7) => N8, A(6) => N9, A(5) => N10, A(4) => N11, 
                           A(3) => N12, A(2) => N13, A(1) => N14, A(0) => N15, 
                           SUM(15) => Y(15), SUM(14) => Y(14), SUM(13) => Y(13)
                           , SUM(12) => Y(12), SUM(11) => Y(11), SUM(10) => 
                           Y(10), SUM(9) => Y(9), SUM(8) => Y(8), SUM(7) => 
                           Y(7), SUM(6) => Y(6), SUM(5) => Y(5), SUM(4) => Y(4)
                           , SUM(3) => Y(3), SUM(2) => Y(2), SUM(1) => Y(1), 
                           SUM(0) => Y(0));
   U2 : INV_X1 port map( A => A(6), ZN => N9);
   U3 : INV_X1 port map( A => A(7), ZN => N8);
   U4 : INV_X1 port map( A => A(8), ZN => N7);
   U5 : INV_X1 port map( A => A(9), ZN => N6);
   U6 : INV_X1 port map( A => A(10), ZN => N5);
   U7 : INV_X1 port map( A => A(11), ZN => N4);
   U8 : INV_X1 port map( A => A(12), ZN => N3);
   U9 : INV_X1 port map( A => A(13), ZN => N2);
   U10 : INV_X1 port map( A => A(0), ZN => N15);
   U11 : INV_X1 port map( A => A(1), ZN => N14);
   U12 : INV_X1 port map( A => A(2), ZN => N13);
   U13 : INV_X1 port map( A => A(3), ZN => N12);
   U14 : INV_X1 port map( A => A(4), ZN => N11);
   U15 : INV_X1 port map( A => A(5), ZN => N10);
   U16 : INV_X1 port map( A => A(14), ZN => N1);
   U17 : INV_X1 port map( A => A(15), ZN => N0);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_1 is

   port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end complementor_N16_1;

architecture SYN_ARCHDATAFLOW of complementor_N16_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component complementor_N16_1_DW01_inc_0
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal N9, N8, N7, N6, N5, N4, N3, N2, N15, N14, N13, N12, N11, N10, N1, N0 
      : std_logic;

begin
   
   add_0_root_add_19_ni : complementor_N16_1_DW01_inc_0 port map( A(15) => N0, 
                           A(14) => N1, A(13) => N2, A(12) => N3, A(11) => N4, 
                           A(10) => N5, A(9) => N6, A(8) => N7, A(7) => N8, 
                           A(6) => N9, A(5) => N10, A(4) => N11, A(3) => N12, 
                           A(2) => N13, A(1) => N14, A(0) => N15, SUM(15) => 
                           Y(15), SUM(14) => Y(14), SUM(13) => Y(13), SUM(12) 
                           => Y(12), SUM(11) => Y(11), SUM(10) => Y(10), SUM(9)
                           => Y(9), SUM(8) => Y(8), SUM(7) => Y(7), SUM(6) => 
                           Y(6), SUM(5) => Y(5), SUM(4) => Y(4), SUM(3) => Y(3)
                           , SUM(2) => Y(2), SUM(1) => Y(1), SUM(0) => Y(0));
   U2 : INV_X1 port map( A => A(6), ZN => N9);
   U3 : INV_X1 port map( A => A(7), ZN => N8);
   U4 : INV_X1 port map( A => A(8), ZN => N7);
   U5 : INV_X1 port map( A => A(9), ZN => N6);
   U6 : INV_X1 port map( A => A(10), ZN => N5);
   U7 : INV_X1 port map( A => A(11), ZN => N4);
   U8 : INV_X1 port map( A => A(12), ZN => N3);
   U9 : INV_X1 port map( A => A(13), ZN => N2);
   U10 : INV_X1 port map( A => A(0), ZN => N15);
   U11 : INV_X1 port map( A => A(1), ZN => N14);
   U12 : INV_X1 port map( A => A(2), ZN => N13);
   U13 : INV_X1 port map( A => A(3), ZN => N12);
   U14 : INV_X1 port map( A => A(4), ZN => N11);
   U15 : INV_X1 port map( A => A(5), ZN => N10);
   U16 : INV_X1 port map( A => A(14), ZN => N1);
   U17 : INV_X1 port map( A => A(15), ZN => N0);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_7 is

   port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector (3 
         downto 0);  SA : out std_logic_vector (15 downto 0));

end shift_pow2_N8_7;

architecture SYN_ARCHBEH of shift_pow2_N8_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_pow2_N8_7_DW02_mult_0_DW02_mult_6
      port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (15 downto 0));
   end component;
   
   signal shift_pow_31_ML_int_4_0_port, shift_pow_31_ML_int_4_1_port, 
      shift_pow_31_ML_int_4_2_port, shift_pow_31_ML_int_4_3_port, 
      shift_pow_31_ML_int_4_4_port, shift_pow_31_ML_int_4_5_port, 
      shift_pow_31_ML_int_4_6_port, shift_pow_31_ML_int_4_7_port, 
      shift_pow_31_ML_int_2_0_port, shift_pow_31_ML_int_2_1_port, n1, n2, n3, 
      n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   n11 <= '0';
   mult_31 : shift_pow2_N8_7_DW02_mult_0_DW02_mult_6 port map( A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), B(7)
                           => shift_pow_31_ML_int_4_7_port, B(6) => 
                           shift_pow_31_ML_int_4_6_port, B(5) => 
                           shift_pow_31_ML_int_4_5_port, B(4) => 
                           shift_pow_31_ML_int_4_4_port, B(3) => 
                           shift_pow_31_ML_int_4_3_port, B(2) => 
                           shift_pow_31_ML_int_4_2_port, B(1) => 
                           shift_pow_31_ML_int_4_1_port, B(0) => 
                           shift_pow_31_ML_int_4_0_port, TC => n11, PRODUCT(15)
                           => SA(15), PRODUCT(14) => SA(14), PRODUCT(13) => 
                           SA(13), PRODUCT(12) => SA(12), PRODUCT(11) => SA(11)
                           , PRODUCT(10) => SA(10), PRODUCT(9) => SA(9), 
                           PRODUCT(8) => SA(8), PRODUCT(7) => SA(7), PRODUCT(6)
                           => SA(6), PRODUCT(5) => SA(5), PRODUCT(4) => SA(4), 
                           PRODUCT(3) => SA(3), PRODUCT(2) => SA(2), PRODUCT(1)
                           => SA(1), PRODUCT(0) => SA(0));
   U3 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_1_port, 
                           ZN => n1);
   U4 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_0_port, 
                           ZN => n2);
   U5 : AND2_X1 port map( A1 => Shift(2), A2 => n6, ZN => n3);
   U7 : AND2_X1 port map( A1 => Shift(2), A2 => n7, ZN => n5);
   U8 : AND2_X1 port map( A1 => Shift(1), A2 => n10, ZN => n6);
   U9 : AND2_X1 port map( A1 => Shift(1), A2 => Shift(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n5, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_7_port);
   U11 : AND2_X1 port map( A1 => n3, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_6_port);
   U12 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_5_port);
   U13 : AND2_X1 port map( A1 => n2, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_4_port);
   U14 : INV_X1 port map( A => Shift(3), ZN => n8);
   U15 : AND2_X1 port map( A1 => n7, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_3_port);
   U16 : AND2_X1 port map( A1 => n6, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_2_port);
   U17 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_1_port, ZN => 
                           shift_pow_31_ML_int_4_1_port);
   U18 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_0_port, ZN => 
                           shift_pow_31_ML_int_4_0_port);
   U19 : NOR2_X1 port map( A1 => Shift(3), A2 => Shift(2), ZN => n9);
   U20 : NOR2_X1 port map( A1 => n10, A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_1_port);
   U21 : NOR2_X1 port map( A1 => Shift(0), A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_0_port);
   U22 : INV_X1 port map( A => Shift(0), ZN => n10);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_6 is

   port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector (3 
         downto 0);  SA : out std_logic_vector (15 downto 0));

end shift_pow2_N8_6;

architecture SYN_ARCHBEH of shift_pow2_N8_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_pow2_N8_6_DW02_mult_0_DW02_mult_5
      port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (15 downto 0));
   end component;
   
   signal shift_pow_31_ML_int_4_0_port, shift_pow_31_ML_int_4_1_port, 
      shift_pow_31_ML_int_4_2_port, shift_pow_31_ML_int_4_3_port, 
      shift_pow_31_ML_int_4_4_port, shift_pow_31_ML_int_4_5_port, 
      shift_pow_31_ML_int_4_6_port, shift_pow_31_ML_int_4_7_port, 
      shift_pow_31_ML_int_2_0_port, shift_pow_31_ML_int_2_1_port, n1, n2, n3, 
      n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   n11 <= '0';
   mult_31 : shift_pow2_N8_6_DW02_mult_0_DW02_mult_5 port map( A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), B(7)
                           => shift_pow_31_ML_int_4_7_port, B(6) => 
                           shift_pow_31_ML_int_4_6_port, B(5) => 
                           shift_pow_31_ML_int_4_5_port, B(4) => 
                           shift_pow_31_ML_int_4_4_port, B(3) => 
                           shift_pow_31_ML_int_4_3_port, B(2) => 
                           shift_pow_31_ML_int_4_2_port, B(1) => 
                           shift_pow_31_ML_int_4_1_port, B(0) => 
                           shift_pow_31_ML_int_4_0_port, TC => n11, PRODUCT(15)
                           => SA(15), PRODUCT(14) => SA(14), PRODUCT(13) => 
                           SA(13), PRODUCT(12) => SA(12), PRODUCT(11) => SA(11)
                           , PRODUCT(10) => SA(10), PRODUCT(9) => SA(9), 
                           PRODUCT(8) => SA(8), PRODUCT(7) => SA(7), PRODUCT(6)
                           => SA(6), PRODUCT(5) => SA(5), PRODUCT(4) => SA(4), 
                           PRODUCT(3) => SA(3), PRODUCT(2) => SA(2), PRODUCT(1)
                           => SA(1), PRODUCT(0) => SA(0));
   U3 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_1_port, 
                           ZN => n1);
   U4 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_0_port, 
                           ZN => n2);
   U5 : AND2_X1 port map( A1 => Shift(2), A2 => n6, ZN => n3);
   U7 : AND2_X1 port map( A1 => Shift(2), A2 => n7, ZN => n5);
   U8 : AND2_X1 port map( A1 => Shift(1), A2 => n10, ZN => n6);
   U9 : AND2_X1 port map( A1 => Shift(1), A2 => Shift(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n5, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_7_port);
   U11 : AND2_X1 port map( A1 => n3, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_6_port);
   U12 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_5_port);
   U13 : AND2_X1 port map( A1 => n2, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_4_port);
   U14 : INV_X1 port map( A => Shift(3), ZN => n8);
   U15 : AND2_X1 port map( A1 => n7, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_3_port);
   U16 : AND2_X1 port map( A1 => n6, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_2_port);
   U17 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_1_port, ZN => 
                           shift_pow_31_ML_int_4_1_port);
   U18 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_0_port, ZN => 
                           shift_pow_31_ML_int_4_0_port);
   U19 : NOR2_X1 port map( A1 => Shift(3), A2 => Shift(2), ZN => n9);
   U20 : NOR2_X1 port map( A1 => n10, A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_1_port);
   U21 : NOR2_X1 port map( A1 => Shift(0), A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_0_port);
   U22 : INV_X1 port map( A => Shift(0), ZN => n10);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_5 is

   port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector (3 
         downto 0);  SA : out std_logic_vector (15 downto 0));

end shift_pow2_N8_5;

architecture SYN_ARCHBEH of shift_pow2_N8_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_pow2_N8_5_DW02_mult_0_DW02_mult_4
      port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (15 downto 0));
   end component;
   
   signal shift_pow_31_ML_int_4_0_port, shift_pow_31_ML_int_4_1_port, 
      shift_pow_31_ML_int_4_2_port, shift_pow_31_ML_int_4_3_port, 
      shift_pow_31_ML_int_4_4_port, shift_pow_31_ML_int_4_5_port, 
      shift_pow_31_ML_int_4_6_port, shift_pow_31_ML_int_4_7_port, 
      shift_pow_31_ML_int_2_0_port, shift_pow_31_ML_int_2_1_port, n1, n2, n3, 
      n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   n11 <= '0';
   mult_31 : shift_pow2_N8_5_DW02_mult_0_DW02_mult_4 port map( A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), B(7)
                           => shift_pow_31_ML_int_4_7_port, B(6) => 
                           shift_pow_31_ML_int_4_6_port, B(5) => 
                           shift_pow_31_ML_int_4_5_port, B(4) => 
                           shift_pow_31_ML_int_4_4_port, B(3) => 
                           shift_pow_31_ML_int_4_3_port, B(2) => 
                           shift_pow_31_ML_int_4_2_port, B(1) => 
                           shift_pow_31_ML_int_4_1_port, B(0) => 
                           shift_pow_31_ML_int_4_0_port, TC => n11, PRODUCT(15)
                           => SA(15), PRODUCT(14) => SA(14), PRODUCT(13) => 
                           SA(13), PRODUCT(12) => SA(12), PRODUCT(11) => SA(11)
                           , PRODUCT(10) => SA(10), PRODUCT(9) => SA(9), 
                           PRODUCT(8) => SA(8), PRODUCT(7) => SA(7), PRODUCT(6)
                           => SA(6), PRODUCT(5) => SA(5), PRODUCT(4) => SA(4), 
                           PRODUCT(3) => SA(3), PRODUCT(2) => SA(2), PRODUCT(1)
                           => SA(1), PRODUCT(0) => SA(0));
   U3 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_1_port, 
                           ZN => n1);
   U4 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_0_port, 
                           ZN => n2);
   U5 : AND2_X1 port map( A1 => Shift(2), A2 => n6, ZN => n3);
   U7 : AND2_X1 port map( A1 => Shift(2), A2 => n7, ZN => n5);
   U8 : AND2_X1 port map( A1 => Shift(1), A2 => n10, ZN => n6);
   U9 : AND2_X1 port map( A1 => Shift(1), A2 => Shift(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n5, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_7_port);
   U11 : AND2_X1 port map( A1 => n3, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_6_port);
   U12 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_5_port);
   U13 : AND2_X1 port map( A1 => n2, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_4_port);
   U14 : INV_X1 port map( A => Shift(3), ZN => n8);
   U15 : AND2_X1 port map( A1 => n7, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_3_port);
   U16 : AND2_X1 port map( A1 => n6, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_2_port);
   U17 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_1_port, ZN => 
                           shift_pow_31_ML_int_4_1_port);
   U18 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_0_port, ZN => 
                           shift_pow_31_ML_int_4_0_port);
   U19 : NOR2_X1 port map( A1 => Shift(3), A2 => Shift(2), ZN => n9);
   U20 : NOR2_X1 port map( A1 => n10, A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_1_port);
   U21 : NOR2_X1 port map( A1 => Shift(0), A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_0_port);
   U22 : INV_X1 port map( A => Shift(0), ZN => n10);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_4 is

   port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector (3 
         downto 0);  SA : out std_logic_vector (15 downto 0));

end shift_pow2_N8_4;

architecture SYN_ARCHBEH of shift_pow2_N8_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_pow2_N8_4_DW02_mult_0_DW02_mult_3
      port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (15 downto 0));
   end component;
   
   signal shift_pow_31_ML_int_4_0_port, shift_pow_31_ML_int_4_1_port, 
      shift_pow_31_ML_int_4_2_port, shift_pow_31_ML_int_4_3_port, 
      shift_pow_31_ML_int_4_4_port, shift_pow_31_ML_int_4_5_port, 
      shift_pow_31_ML_int_4_6_port, shift_pow_31_ML_int_4_7_port, 
      shift_pow_31_ML_int_2_0_port, shift_pow_31_ML_int_2_1_port, n1, n2, n3, 
      n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   n11 <= '0';
   mult_31 : shift_pow2_N8_4_DW02_mult_0_DW02_mult_3 port map( A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), B(7)
                           => shift_pow_31_ML_int_4_7_port, B(6) => 
                           shift_pow_31_ML_int_4_6_port, B(5) => 
                           shift_pow_31_ML_int_4_5_port, B(4) => 
                           shift_pow_31_ML_int_4_4_port, B(3) => 
                           shift_pow_31_ML_int_4_3_port, B(2) => 
                           shift_pow_31_ML_int_4_2_port, B(1) => 
                           shift_pow_31_ML_int_4_1_port, B(0) => 
                           shift_pow_31_ML_int_4_0_port, TC => n11, PRODUCT(15)
                           => SA(15), PRODUCT(14) => SA(14), PRODUCT(13) => 
                           SA(13), PRODUCT(12) => SA(12), PRODUCT(11) => SA(11)
                           , PRODUCT(10) => SA(10), PRODUCT(9) => SA(9), 
                           PRODUCT(8) => SA(8), PRODUCT(7) => SA(7), PRODUCT(6)
                           => SA(6), PRODUCT(5) => SA(5), PRODUCT(4) => SA(4), 
                           PRODUCT(3) => SA(3), PRODUCT(2) => SA(2), PRODUCT(1)
                           => SA(1), PRODUCT(0) => SA(0));
   U3 : AND2_X1 port map( A1 => Shift(2), A2 => n6, ZN => n1);
   U4 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_1_port, 
                           ZN => n2);
   U5 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_0_port, 
                           ZN => n3);
   U7 : AND2_X1 port map( A1 => Shift(2), A2 => n7, ZN => n5);
   U8 : AND2_X1 port map( A1 => Shift(1), A2 => n10, ZN => n6);
   U9 : AND2_X1 port map( A1 => Shift(1), A2 => Shift(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n5, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_7_port);
   U11 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_6_port);
   U12 : AND2_X1 port map( A1 => n2, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_5_port);
   U13 : AND2_X1 port map( A1 => n3, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_4_port);
   U14 : INV_X1 port map( A => Shift(3), ZN => n8);
   U15 : AND2_X1 port map( A1 => n7, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_3_port);
   U16 : AND2_X1 port map( A1 => n6, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_2_port);
   U17 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_1_port, ZN => 
                           shift_pow_31_ML_int_4_1_port);
   U18 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_0_port, ZN => 
                           shift_pow_31_ML_int_4_0_port);
   U19 : NOR2_X1 port map( A1 => Shift(3), A2 => Shift(2), ZN => n9);
   U20 : NOR2_X1 port map( A1 => n10, A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_1_port);
   U21 : NOR2_X1 port map( A1 => Shift(0), A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_0_port);
   U22 : INV_X1 port map( A => Shift(0), ZN => n10);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_3 is

   port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector (3 
         downto 0);  SA : out std_logic_vector (15 downto 0));

end shift_pow2_N8_3;

architecture SYN_ARCHBEH of shift_pow2_N8_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_pow2_N8_3_DW02_mult_0_DW02_mult_2
      port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (15 downto 0));
   end component;
   
   signal shift_pow_31_ML_int_4_0_port, shift_pow_31_ML_int_4_1_port, 
      shift_pow_31_ML_int_4_2_port, shift_pow_31_ML_int_4_3_port, 
      shift_pow_31_ML_int_4_4_port, shift_pow_31_ML_int_4_5_port, 
      shift_pow_31_ML_int_4_6_port, shift_pow_31_ML_int_4_7_port, 
      shift_pow_31_ML_int_2_0_port, shift_pow_31_ML_int_2_1_port, n1, n2, n3, 
      n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   n11 <= '0';
   mult_31 : shift_pow2_N8_3_DW02_mult_0_DW02_mult_2 port map( A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), B(7)
                           => shift_pow_31_ML_int_4_7_port, B(6) => 
                           shift_pow_31_ML_int_4_6_port, B(5) => 
                           shift_pow_31_ML_int_4_5_port, B(4) => 
                           shift_pow_31_ML_int_4_4_port, B(3) => 
                           shift_pow_31_ML_int_4_3_port, B(2) => 
                           shift_pow_31_ML_int_4_2_port, B(1) => 
                           shift_pow_31_ML_int_4_1_port, B(0) => 
                           shift_pow_31_ML_int_4_0_port, TC => n11, PRODUCT(15)
                           => SA(15), PRODUCT(14) => SA(14), PRODUCT(13) => 
                           SA(13), PRODUCT(12) => SA(12), PRODUCT(11) => SA(11)
                           , PRODUCT(10) => SA(10), PRODUCT(9) => SA(9), 
                           PRODUCT(8) => SA(8), PRODUCT(7) => SA(7), PRODUCT(6)
                           => SA(6), PRODUCT(5) => SA(5), PRODUCT(4) => SA(4), 
                           PRODUCT(3) => SA(3), PRODUCT(2) => SA(2), PRODUCT(1)
                           => SA(1), PRODUCT(0) => SA(0));
   U3 : AND2_X1 port map( A1 => Shift(2), A2 => n6, ZN => n1);
   U4 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_1_port, 
                           ZN => n2);
   U5 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_0_port, 
                           ZN => n3);
   U7 : AND2_X1 port map( A1 => Shift(2), A2 => n7, ZN => n5);
   U8 : AND2_X1 port map( A1 => Shift(1), A2 => n10, ZN => n6);
   U9 : AND2_X1 port map( A1 => Shift(1), A2 => Shift(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n5, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_7_port);
   U11 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_6_port);
   U12 : AND2_X1 port map( A1 => n2, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_5_port);
   U13 : AND2_X1 port map( A1 => n3, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_4_port);
   U14 : INV_X1 port map( A => Shift(3), ZN => n8);
   U15 : AND2_X1 port map( A1 => n7, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_3_port);
   U16 : AND2_X1 port map( A1 => n6, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_2_port);
   U17 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_1_port, ZN => 
                           shift_pow_31_ML_int_4_1_port);
   U18 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_0_port, ZN => 
                           shift_pow_31_ML_int_4_0_port);
   U19 : NOR2_X1 port map( A1 => Shift(3), A2 => Shift(2), ZN => n9);
   U20 : NOR2_X1 port map( A1 => n10, A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_1_port);
   U21 : NOR2_X1 port map( A1 => Shift(0), A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_0_port);
   U22 : INV_X1 port map( A => Shift(0), ZN => n10);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_2 is

   port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector (3 
         downto 0);  SA : out std_logic_vector (15 downto 0));

end shift_pow2_N8_2;

architecture SYN_ARCHBEH of shift_pow2_N8_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_pow2_N8_2_DW02_mult_0_DW02_mult_1
      port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (15 downto 0));
   end component;
   
   signal shift_pow_31_ML_int_4_0_port, shift_pow_31_ML_int_4_1_port, 
      shift_pow_31_ML_int_4_2_port, shift_pow_31_ML_int_4_3_port, 
      shift_pow_31_ML_int_4_4_port, shift_pow_31_ML_int_4_5_port, 
      shift_pow_31_ML_int_4_6_port, shift_pow_31_ML_int_4_7_port, 
      shift_pow_31_ML_int_2_0_port, shift_pow_31_ML_int_2_1_port, n1, n2, n3, 
      n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   n11 <= '0';
   mult_31 : shift_pow2_N8_2_DW02_mult_0_DW02_mult_1 port map( A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), B(7)
                           => shift_pow_31_ML_int_4_7_port, B(6) => 
                           shift_pow_31_ML_int_4_6_port, B(5) => 
                           shift_pow_31_ML_int_4_5_port, B(4) => 
                           shift_pow_31_ML_int_4_4_port, B(3) => 
                           shift_pow_31_ML_int_4_3_port, B(2) => 
                           shift_pow_31_ML_int_4_2_port, B(1) => 
                           shift_pow_31_ML_int_4_1_port, B(0) => 
                           shift_pow_31_ML_int_4_0_port, TC => n11, PRODUCT(15)
                           => SA(15), PRODUCT(14) => SA(14), PRODUCT(13) => 
                           SA(13), PRODUCT(12) => SA(12), PRODUCT(11) => SA(11)
                           , PRODUCT(10) => SA(10), PRODUCT(9) => SA(9), 
                           PRODUCT(8) => SA(8), PRODUCT(7) => SA(7), PRODUCT(6)
                           => SA(6), PRODUCT(5) => SA(5), PRODUCT(4) => SA(4), 
                           PRODUCT(3) => SA(3), PRODUCT(2) => SA(2), PRODUCT(1)
                           => SA(1), PRODUCT(0) => SA(0));
   U3 : AND2_X1 port map( A1 => Shift(2), A2 => n6, ZN => n1);
   U4 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_1_port, 
                           ZN => n2);
   U5 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_0_port, 
                           ZN => n3);
   U7 : AND2_X1 port map( A1 => Shift(2), A2 => n7, ZN => n5);
   U8 : AND2_X1 port map( A1 => Shift(1), A2 => n10, ZN => n6);
   U9 : AND2_X1 port map( A1 => Shift(1), A2 => Shift(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n5, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_7_port);
   U11 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_6_port);
   U12 : AND2_X1 port map( A1 => n2, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_5_port);
   U13 : AND2_X1 port map( A1 => n3, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_4_port);
   U14 : INV_X1 port map( A => Shift(3), ZN => n8);
   U15 : AND2_X1 port map( A1 => n7, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_3_port);
   U16 : AND2_X1 port map( A1 => n6, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_2_port);
   U17 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_1_port, ZN => 
                           shift_pow_31_ML_int_4_1_port);
   U18 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_0_port, ZN => 
                           shift_pow_31_ML_int_4_0_port);
   U19 : NOR2_X1 port map( A1 => Shift(3), A2 => Shift(2), ZN => n9);
   U20 : NOR2_X1 port map( A1 => n10, A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_1_port);
   U21 : NOR2_X1 port map( A1 => Shift(0), A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_0_port);
   U22 : INV_X1 port map( A => Shift(0), ZN => n10);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_1 is

   port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector (3 
         downto 0);  SA : out std_logic_vector (15 downto 0));

end shift_pow2_N8_1;

architecture SYN_ARCHBEH of shift_pow2_N8_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_pow2_N8_1_DW02_mult_0
      port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (15 downto 0));
   end component;
   
   signal shift_pow_31_ML_int_4_0_port, shift_pow_31_ML_int_4_1_port, 
      shift_pow_31_ML_int_4_2_port, shift_pow_31_ML_int_4_3_port, 
      shift_pow_31_ML_int_4_4_port, shift_pow_31_ML_int_4_5_port, 
      shift_pow_31_ML_int_4_6_port, shift_pow_31_ML_int_4_7_port, 
      shift_pow_31_ML_int_2_0_port, shift_pow_31_ML_int_2_1_port, n1, n2, n3, 
      n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   n11 <= '0';
   mult_31 : shift_pow2_N8_1_DW02_mult_0 port map( A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(7) => 
                           shift_pow_31_ML_int_4_7_port, B(6) => 
                           shift_pow_31_ML_int_4_6_port, B(5) => 
                           shift_pow_31_ML_int_4_5_port, B(4) => 
                           shift_pow_31_ML_int_4_4_port, B(3) => 
                           shift_pow_31_ML_int_4_3_port, B(2) => 
                           shift_pow_31_ML_int_4_2_port, B(1) => 
                           shift_pow_31_ML_int_4_1_port, B(0) => 
                           shift_pow_31_ML_int_4_0_port, TC => n11, PRODUCT(15)
                           => SA(15), PRODUCT(14) => SA(14), PRODUCT(13) => 
                           SA(13), PRODUCT(12) => SA(12), PRODUCT(11) => SA(11)
                           , PRODUCT(10) => SA(10), PRODUCT(9) => SA(9), 
                           PRODUCT(8) => SA(8), PRODUCT(7) => SA(7), PRODUCT(6)
                           => SA(6), PRODUCT(5) => SA(5), PRODUCT(4) => SA(4), 
                           PRODUCT(3) => SA(3), PRODUCT(2) => SA(2), PRODUCT(1)
                           => SA(1), PRODUCT(0) => SA(0));
   U3 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_1_port, 
                           ZN => n1);
   U4 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_0_port, 
                           ZN => n2);
   U5 : AND2_X1 port map( A1 => Shift(2), A2 => n6, ZN => n3);
   U7 : AND2_X1 port map( A1 => Shift(2), A2 => n7, ZN => n5);
   U8 : AND2_X1 port map( A1 => Shift(1), A2 => n10, ZN => n6);
   U9 : AND2_X1 port map( A1 => Shift(1), A2 => Shift(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n5, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_7_port);
   U11 : AND2_X1 port map( A1 => n3, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_6_port);
   U12 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_5_port);
   U13 : AND2_X1 port map( A1 => n2, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_4_port);
   U14 : INV_X1 port map( A => Shift(3), ZN => n8);
   U15 : AND2_X1 port map( A1 => n7, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_3_port);
   U16 : AND2_X1 port map( A1 => n6, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_2_port);
   U17 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_1_port, ZN => 
                           shift_pow_31_ML_int_4_1_port);
   U18 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_0_port, ZN => 
                           shift_pow_31_ML_int_4_0_port);
   U19 : NOR2_X1 port map( A1 => Shift(3), A2 => Shift(2), ZN => n9);
   U20 : NOR2_X1 port map( A1 => n10, A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_1_port);
   U21 : NOR2_X1 port map( A1 => Shift(0), A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_0_port);
   U22 : INV_X1 port map( A => Shift(0), ZN => n10);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity FA_1920 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1920;

architecture SYN_ARCHBEH of FA_1920 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n1);
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N4_240 is

   port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (3 downto 0));

end muxN1_N4_240;

architecture SYN_ARCHSTRUCT of muxN1_N4_240 is

   component mux21_8173
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8174
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8175
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8176
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   mux21_g_0 : mux21_8176 port map( A => A(0), B => B(0), S => S, Y => Y(0));
   mux21_g_1 : mux21_8175 port map( A => A(1), B => B(1), S => S, Y => Y(1));
   mux21_g_2 : mux21_8174 port map( A => A(2), B => B(2), S => S, Y => Y(2));
   mux21_g_3 : mux21_8173 port map( A => A(3), B => B(3), S => S, Y => Y(3));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity RCA_N4_480 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_N4_480;

architecture SYN_ARCHSTRUCT of RCA_N4_480 is

   component FA_2013
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2014
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2015
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1920
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_1920 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_2015 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_2014 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_2013 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => Co);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_block_945 is

   port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : out
         std_logic);

end pg_block_945;

architecture SYN_ARCHDATAFLOW of pg_block_945 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);
   U3 : AND2_X1 port map( A1 => P_kmin1_j, A2 => P_i_k, ZN => P_i_j);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity g_block_255 is

   port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);

end g_block_255;

architecture SYN_ARCHDATAFLOW of g_block_255 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_i_j);
   U2 : AOI21_X1 port map( B1 => P_i_k, B2 => G_kmin1_j, A => G_i_k, ZN => n1);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity nd2_24384 is

   port( A, B : in std_logic;  Y : out std_logic);

end nd2_24384;

architecture SYN_ARCHBEH of nd2_24384 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity iv_8128 is

   port( A : in std_logic;  Y : out std_logic);

end iv_8128;

architecture SYN_ARCHSTRUCT of iv_8128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_select_block_N4_240 is

   port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : out
         std_logic_vector (3 downto 0));

end carry_select_block_N4_240;

architecture SYN_ARCHSTRUCT of carry_select_block_N4_240 is

   component muxN1_N4_240
      port( A, B : in std_logic_vector (3 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_N4_503
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_N4_480
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S1_3_port, S1_2_port, S1_1_port, 
      S1_0_port, S2_3_port, S2_2_port, S2_1_port, S2_0_port, n_1120, n_1121 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_N4_480 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => S1_3_port
                           , S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1120);
   RCA2 : RCA_N4_503 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => S2_3_port
                           , S(2) => S2_2_port, S(1) => S2_1_port, S(0) => 
                           S2_0_port, Co => n_1121);
   MUX : muxN1_N4_240 port map( A(3) => S2_3_port, A(2) => S2_2_port, A(1) => 
                           S2_1_port, A(0) => S2_0_port, B(3) => S1_3_port, 
                           B(2) => S1_2_port, B(1) => S1_1_port, B(0) => 
                           S1_0_port, S => Cin, Y(3) => S(3), Y(2) => S(2), 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_generator_sparse_tree_N16_carry_range4_0 is

   port( P, G : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C : 
         out std_logic_vector (4 downto 0));

end carry_generator_sparse_tree_N16_carry_range4_0;

architecture SYN_ARCHSTRUCT of carry_generator_sparse_tree_N16_carry_range4_0 
   is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component g_block_266
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component g_block_267
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_968
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_268
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_969
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_970
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_971
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_269
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   component pg_block_972
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_973
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_974
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_975
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_976
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_977
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component pg_block_945
      port( G_i_k, G_kmin1_j, P_i_k, P_kmin1_j : in std_logic;  P_i_j, G_i_j : 
            out std_logic);
   end component;
   
   component g_block_255
      port( G_i_k, G_kmin1_j, P_i_k : in std_logic;  G_i_j : out std_logic);
   end component;
   
   signal C_4_port, C_3_port, C_2_port, C_1_port, Gmat_16_15_port, 
      Gmat_16_13_port, Gmat_16_9_port, Gmat_14_13_port, Gmat_12_11_port, 
      Gmat_12_9_port, Gmat_10_9_port, Gmat_8_7_port, Gmat_8_5_port, 
      Gmat_6_5_port, Gmat_4_3_port, Gmat_2_1_port, Pmat_16_15_port, 
      Pmat_16_13_port, Pmat_16_9_port, Pmat_14_13_port, Pmat_12_11_port, 
      Pmat_12_9_port, Pmat_10_9_port, Pmat_8_7_port, Pmat_8_5_port, 
      Pmat_6_5_port, Pmat_4_3_port, n1, n2 : std_logic;

begin
   C <= ( C_4_port, C_3_port, C_2_port, C_1_port, Cin );
   
   first_G_1_2 : g_block_255 port map( G_i_k => G(1), G_kmin1_j => n2, P_i_k =>
                           P(1), G_i_j => Gmat_2_1_port);
   FRST_PG_1_4 : pg_block_945 port map( G_i_k => G(3), G_kmin1_j => G(2), P_i_k
                           => P(3), P_kmin1_j => P(2), P_i_j => Pmat_4_3_port, 
                           G_i_j => Gmat_4_3_port);
   FRST_PG_1_6 : pg_block_977 port map( G_i_k => G(5), G_kmin1_j => G(4), P_i_k
                           => P(5), P_kmin1_j => P(4), P_i_j => Pmat_6_5_port, 
                           G_i_j => Gmat_6_5_port);
   FRST_PG_1_8 : pg_block_976 port map( G_i_k => G(7), G_kmin1_j => G(6), P_i_k
                           => P(7), P_kmin1_j => P(6), P_i_j => Pmat_8_7_port, 
                           G_i_j => Gmat_8_7_port);
   FRST_PG_1_10 : pg_block_975 port map( G_i_k => G(9), G_kmin1_j => G(8), 
                           P_i_k => P(9), P_kmin1_j => P(8), P_i_j => 
                           Pmat_10_9_port, G_i_j => Gmat_10_9_port);
   FRST_PG_1_12 : pg_block_974 port map( G_i_k => G(11), G_kmin1_j => G(10), 
                           P_i_k => P(11), P_kmin1_j => P(10), P_i_j => 
                           Pmat_12_11_port, G_i_j => Gmat_12_11_port);
   FRST_PG_1_14 : pg_block_973 port map( G_i_k => G(13), G_kmin1_j => G(12), 
                           P_i_k => P(13), P_kmin1_j => P(12), P_i_j => 
                           Pmat_14_13_port, G_i_j => Gmat_14_13_port);
   FRST_PG_1_16 : pg_block_972 port map( G_i_k => G(15), G_kmin1_j => G(14), 
                           P_i_k => P(15), P_kmin1_j => P(14), P_i_j => 
                           Pmat_16_15_port, G_i_j => Gmat_16_15_port);
   first_G_2_4 : g_block_269 port map( G_i_k => Gmat_4_3_port, G_kmin1_j => 
                           Gmat_2_1_port, P_i_k => Pmat_4_3_port, G_i_j => 
                           C_1_port);
   FRST_PG_2_8 : pg_block_971 port map( G_i_k => Gmat_8_7_port, G_kmin1_j => 
                           Gmat_6_5_port, P_i_k => Pmat_8_7_port, P_kmin1_j => 
                           Pmat_6_5_port, P_i_j => Pmat_8_5_port, G_i_j => 
                           Gmat_8_5_port);
   FRST_PG_2_12 : pg_block_970 port map( G_i_k => Gmat_12_11_port, G_kmin1_j =>
                           Gmat_10_9_port, P_i_k => Pmat_12_11_port, P_kmin1_j 
                           => Pmat_10_9_port, P_i_j => Pmat_12_9_port, G_i_j =>
                           Gmat_12_9_port);
   FRST_PG_2_16 : pg_block_969 port map( G_i_k => Gmat_16_15_port, G_kmin1_j =>
                           Gmat_14_13_port, P_i_k => Pmat_16_15_port, P_kmin1_j
                           => Pmat_14_13_port, P_i_j => Pmat_16_13_port, G_i_j 
                           => Gmat_16_13_port);
   G_L2_0_4_8 : g_block_268 port map( G_i_k => Gmat_8_5_port, G_kmin1_j => 
                           C_1_port, P_i_k => Pmat_8_5_port, G_i_j => C_2_port)
                           ;
   PG_L2_0_12_16 : pg_block_968 port map( G_i_k => Gmat_16_13_port, G_kmin1_j 
                           => Gmat_12_9_port, P_i_k => Pmat_16_13_port, 
                           P_kmin1_j => Pmat_12_9_port, P_i_j => Pmat_16_9_port
                           , G_i_j => Gmat_16_9_port);
   G_L2_1_8_12 : g_block_267 port map( G_i_k => Gmat_12_9_port, G_kmin1_j => 
                           C_2_port, P_i_k => Pmat_12_9_port, G_i_j => C_3_port
                           );
   G_L2_1_8_16 : g_block_266 port map( G_i_k => Gmat_16_9_port, G_kmin1_j => 
                           C_2_port, P_i_k => Pmat_16_9_port, G_i_j => C_4_port
                           );
   U1 : INV_X1 port map( A => n1, ZN => n2);
   U2 : AOI21_X1 port map( B1 => P(0), B2 => Cin, A => G(0), ZN => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity pg_network_N16_0 is

   port( A, B : in std_logic_vector (15 downto 0);  P, G : out std_logic_vector
         (15 downto 0));

end pg_network_N16_0;

architecture SYN_ARCHDATAFLOW of pg_network_N16_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B(9), B => A(9), Z => P(9));
   U2 : XOR2_X1 port map( A => B(8), B => A(8), Z => P(8));
   U3 : XOR2_X1 port map( A => B(7), B => A(7), Z => P(7));
   U4 : XOR2_X1 port map( A => B(6), B => A(6), Z => P(6));
   U5 : XOR2_X1 port map( A => B(5), B => A(5), Z => P(5));
   U6 : XOR2_X1 port map( A => B(4), B => A(4), Z => P(4));
   U7 : XOR2_X1 port map( A => B(3), B => A(3), Z => P(3));
   U8 : XOR2_X1 port map( A => B(2), B => A(2), Z => P(2));
   U9 : XOR2_X1 port map( A => B(1), B => A(1), Z => P(1));
   U10 : XOR2_X1 port map( A => B(15), B => A(15), Z => P(15));
   U11 : XOR2_X1 port map( A => B(14), B => A(14), Z => P(14));
   U12 : XOR2_X1 port map( A => B(13), B => A(13), Z => P(13));
   U13 : XOR2_X1 port map( A => B(12), B => A(12), Z => P(12));
   U14 : XOR2_X1 port map( A => B(11), B => A(11), Z => P(11));
   U15 : XOR2_X1 port map( A => B(10), B => A(10), Z => P(10));
   U16 : XOR2_X1 port map( A => B(0), B => A(0), Z => P(0));
   U17 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => G(9));
   U18 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => G(8));
   U19 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => G(7));
   U20 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => G(6));
   U21 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => G(5));
   U22 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => G(4));
   U23 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => G(3));
   U24 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => G(2));
   U25 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => G(1));
   U26 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => G(15));
   U27 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => G(14));
   U28 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => G(13));
   U29 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => G(12));
   U30 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => G(11));
   U31 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => G(10));
   U32 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => G(0));

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux21_8128 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end mux21_8128;

architecture SYN_ARCHSTRUCT of mux21_8128 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nd2_25870
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_25871
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component nd2_24384
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component iv_8128
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal n_S, s1, s2, n1 : std_logic;

begin
   
   NOT1 : iv_8128 port map( A => n1, Y => n_S);
   NAND1 : nd2_24384 port map( A => A, B => n1, Y => s1);
   NAND2 : nd2_25871 port map( A => B, B => n_S, Y => s2);
   NAND3 : nd2_25870 port map( A => s1, B => s2, Y => Y);
   U1 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity sum_generator_N16_Nbit_blocks4_0 is

   port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  Carry 
         : in std_logic_vector (3 downto 0);  S : out std_logic_vector (15 
         downto 0);  Cout : out std_logic);

end sum_generator_N16_Nbit_blocks4_0;

architecture SYN_ARCHSTRUCT of sum_generator_N16_Nbit_blocks4_0 is

   component carry_select_block_N4_249
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_250
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_251
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_N4_240
      port( Cin : in std_logic;  A, B : in std_logic_vector (3 downto 0);  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   Cout <= Carry(3);
   
   CSB_1 : carry_select_block_N4_240 port map( Cin => Cin, A(3) => A(3), A(2) 
                           => A(2), A(1) => A(1), A(0) => A(0), B(3) => B(3), 
                           B(2) => B(2), B(1) => B(1), B(0) => B(0), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   CSB_2 : carry_select_block_N4_251 port map( Cin => Carry(0), A(3) => A(7), 
                           A(2) => A(6), A(1) => A(5), A(0) => A(4), B(3) => 
                           B(7), B(2) => B(6), B(1) => B(5), B(0) => B(4), S(3)
                           => S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   CSB_3 : carry_select_block_N4_250 port map( Cin => Carry(1), A(3) => A(11), 
                           A(2) => A(10), A(1) => A(9), A(0) => A(8), B(3) => 
                           B(11), B(2) => B(10), B(1) => B(9), B(0) => B(8), 
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   CSB_4 : carry_select_block_N4_249 port map( Cin => Carry(2), A(3) => A(15), 
                           A(2) => A(14), A(1) => A(13), A(0) => A(12), B(3) =>
                           B(15), B(2) => B(14), B(1) => B(13), B(0) => B(12), 
                           S(3) => S(15), S(2) => S(14), S(1) => S(13), S(0) =>
                           S(12));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity carry_generator_N16_carry_range4_0 is

   port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C : 
         out std_logic_vector (4 downto 0));

end carry_generator_N16_carry_range4_0;

architecture SYN_ARCHSTRUCT of carry_generator_N16_carry_range4_0 is

   component carry_generator_sparse_tree_N16_carry_range4_0
      port( P, G : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C :
            out std_logic_vector (4 downto 0));
   end component;
   
   component pg_network_N16_0
      port( A, B : in std_logic_vector (15 downto 0);  P, G : out 
            std_logic_vector (15 downto 0));
   end component;
   
   signal P_15_port, P_14_port, P_13_port, P_12_port, P_11_port, P_10_port, 
      P_9_port, P_8_port, P_7_port, P_6_port, P_5_port, P_4_port, P_3_port, 
      P_2_port, P_1_port, P_0_port, G_15_port, G_14_port, G_13_port, G_12_port,
      G_11_port, G_10_port, G_9_port, G_8_port, G_7_port, G_6_port, G_5_port, 
      G_4_port, G_3_port, G_2_port, G_1_port, G_0_port : std_logic;

begin
   
   PG_NET : pg_network_N16_0 port map( A(15) => A(15), A(14) => A(14), A(13) =>
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), P(15) => P_15_port
                           , P(14) => P_14_port, P(13) => P_13_port, P(12) => 
                           P_12_port, P(11) => P_11_port, P(10) => P_10_port, 
                           P(9) => P_9_port, P(8) => P_8_port, P(7) => P_7_port
                           , P(6) => P_6_port, P(5) => P_5_port, P(4) => 
                           P_4_port, P(3) => P_3_port, P(2) => P_2_port, P(1) 
                           => P_1_port, P(0) => P_0_port, G(15) => G_15_port, 
                           G(14) => G_14_port, G(13) => G_13_port, G(12) => 
                           G_12_port, G(11) => G_11_port, G(10) => G_10_port, 
                           G(9) => G_9_port, G(8) => G_8_port, G(7) => G_7_port
                           , G(6) => G_6_port, G(5) => G_5_port, G(4) => 
                           G_4_port, G(3) => G_3_port, G(2) => G_2_port, G(1) 
                           => G_1_port, G(0) => G_0_port);
   CG : carry_generator_sparse_tree_N16_carry_range4_0 port map( P(15) => 
                           P_15_port, P(14) => P_14_port, P(13) => P_13_port, 
                           P(12) => P_12_port, P(11) => P_11_port, P(10) => 
                           P_10_port, P(9) => P_9_port, P(8) => P_8_port, P(7) 
                           => P_7_port, P(6) => P_6_port, P(5) => P_5_port, 
                           P(4) => P_4_port, P(3) => P_3_port, P(2) => P_2_port
                           , P(1) => P_1_port, P(0) => P_0_port, G(15) => 
                           G_15_port, G(14) => G_14_port, G(13) => G_13_port, 
                           G(12) => G_12_port, G(11) => G_11_port, G(10) => 
                           G_10_port, G(9) => G_9_port, G(8) => G_8_port, G(7) 
                           => G_7_port, G(6) => G_6_port, G(5) => G_5_port, 
                           G(4) => G_4_port, G(3) => G_3_port, G(2) => G_2_port
                           , G(1) => G_1_port, G(0) => G_0_port, Cin => Cin, 
                           C(4) => C(4), C(3) => C(3), C(2) => C(2), C(1) => 
                           C(1), C(0) => C(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity muxN1_N16_0 is

   port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (15 downto 0));

end muxN1_N16_0;

architecture SYN_ARCHSTRUCT of muxN1_N16_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_8609
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8610
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8611
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8612
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8613
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8614
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8615
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8616
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8617
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8618
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8619
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8620
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8621
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8622
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8623
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component mux21_8128
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   mux21_g_0 : mux21_8128 port map( A => A(0), B => B(0), S => n3, Y => Y(0));
   mux21_g_1 : mux21_8623 port map( A => A(1), B => B(1), S => n2, Y => Y(1));
   mux21_g_2 : mux21_8622 port map( A => A(2), B => B(2), S => n2, Y => Y(2));
   mux21_g_3 : mux21_8621 port map( A => A(3), B => B(3), S => n2, Y => Y(3));
   mux21_g_4 : mux21_8620 port map( A => A(4), B => B(4), S => n2, Y => Y(4));
   mux21_g_5 : mux21_8619 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   mux21_g_6 : mux21_8618 port map( A => A(6), B => B(6), S => n2, Y => Y(6));
   mux21_g_7 : mux21_8617 port map( A => A(7), B => B(7), S => n2, Y => Y(7));
   mux21_g_8 : mux21_8616 port map( A => A(8), B => B(8), S => n2, Y => Y(8));
   mux21_g_9 : mux21_8615 port map( A => A(9), B => B(9), S => n2, Y => Y(9));
   mux21_g_10 : mux21_8614 port map( A => A(10), B => B(10), S => n2, Y => 
                           Y(10));
   mux21_g_11 : mux21_8613 port map( A => A(11), B => B(11), S => n2, Y => 
                           Y(11));
   mux21_g_12 : mux21_8612 port map( A => A(12), B => B(12), S => n2, Y => 
                           Y(12));
   mux21_g_13 : mux21_8611 port map( A => A(13), B => B(13), S => n3, Y => 
                           Y(13));
   mux21_g_14 : mux21_8610 port map( A => A(14), B => B(14), S => n3, Y => 
                           Y(14));
   mux21_g_15 : mux21_8609 port map( A => A(15), B => B(15), S => n3, Y => 
                           Y(15));
   U1 : BUF_X1 port map( A => n1, Z => n2);
   U2 : BUF_X1 port map( A => n1, Z => n3);
   U3 : BUF_X1 port map( A => S, Z => n1);

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity booth_encoder_block_16 is

   port( Bi : in std_logic_vector (2 downto 0);  So : out std_logic_vector (2 
         downto 0));

end booth_encoder_block_16;

architecture SYN_DATAFLOW of booth_encoder_block_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U3 : INV_X4 port map( A => Bi(1), ZN => So(1));
   U4 : INV_X2 port map( A => Bi(2), ZN => So(2));
   U5 : INV_X1 port map( A => Bi(0), ZN => So(0));

end SYN_DATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity P4_adder_N16_Nbit_blocks4_0 is

   port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (15 downto 0);  Cout : out std_logic);

end P4_adder_N16_Nbit_blocks4_0;

architecture SYN_STRUCT of P4_adder_N16_Nbit_blocks4_0 is

   component sum_generator_N16_Nbit_blocks4_0
      port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  
            Carry : in std_logic_vector (3 downto 0);  S : out std_logic_vector
            (15 downto 0);  Cout : out std_logic);
   end component;
   
   component carry_generator_N16_carry_range4_0
      port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  C :
            out std_logic_vector (4 downto 0));
   end component;
   
   signal Carries_4_port, Carries_3_port, Carries_2_port, Carries_1_port, 
      n_1122 : std_logic;

begin
   
   CG : carry_generator_N16_carry_range4_0 port map( A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), Cin 
                           => Cin, C(4) => Carries_4_port, C(3) => 
                           Carries_3_port, C(2) => Carries_2_port, C(1) => 
                           Carries_1_port, C(0) => n_1122);
   SG : sum_generator_N16_Nbit_blocks4_0 port map( A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), Cin 
                           => Cin, Carry(3) => Carries_4_port, Carry(2) => 
                           Carries_3_port, Carry(1) => Carries_2_port, Carry(0)
                           => Carries_1_port, S(15) => S(15), S(14) => S(14), 
                           S(13) => S(13), S(12) => S(12), S(11) => S(11), 
                           S(10) => S(10), S(9) => S(9), S(8) => S(8), S(7) => 
                           S(7), S(6) => S(6), S(5) => S(5), S(4) => S(4), S(3)
                           => S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0), 
                           Cout => Cout);

end SYN_STRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity mux_8to1_N16_0 is

   port( A1, A2, A3, A4, A5, A6, A7, A8 : in std_logic_vector (15 downto 0);  S
         : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end mux_8to1_N16_0;

architecture SYN_ARCHSTRUCT of mux_8to1_N16_0 is

   component muxN1_N16_22
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_23
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_24
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_25
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_26
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_27
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   component muxN1_N16_0
      port( A, B : in std_logic_vector (15 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (15 downto 0));
   end component;
   
   signal out1_15_port, out1_14_port, out1_13_port, out1_12_port, out1_11_port,
      out1_10_port, out1_9_port, out1_8_port, out1_7_port, out1_6_port, 
      out1_5_port, out1_4_port, out1_3_port, out1_2_port, out1_1_port, 
      out1_0_port, out2_15_port, out2_14_port, out2_13_port, out2_12_port, 
      out2_11_port, out2_10_port, out2_9_port, out2_8_port, out2_7_port, 
      out2_6_port, out2_5_port, out2_4_port, out2_3_port, out2_2_port, 
      out2_1_port, out2_0_port, out3_15_port, out3_14_port, out3_13_port, 
      out3_12_port, out3_11_port, out3_10_port, out3_9_port, out3_8_port, 
      out3_7_port, out3_6_port, out3_5_port, out3_4_port, out3_3_port, 
      out3_2_port, out3_1_port, out3_0_port, out4_15_port, out4_14_port, 
      out4_13_port, out4_12_port, out4_11_port, out4_10_port, out4_9_port, 
      out4_8_port, out4_7_port, out4_6_port, out4_5_port, out4_4_port, 
      out4_3_port, out4_2_port, out4_1_port, out4_0_port, out5_15_port, 
      out5_14_port, out5_13_port, out5_12_port, out5_11_port, out5_10_port, 
      out5_9_port, out5_8_port, out5_7_port, out5_6_port, out5_5_port, 
      out5_4_port, out5_3_port, out5_2_port, out5_1_port, out5_0_port, 
      out6_15_port, out6_14_port, out6_13_port, out6_12_port, out6_11_port, 
      out6_10_port, out6_9_port, out6_8_port, out6_7_port, out6_6_port, 
      out6_5_port, out6_4_port, out6_3_port, out6_2_port, out6_1_port, 
      out6_0_port : std_logic;

begin
   
   MUX1 : muxN1_N16_0 port map( A(15) => A1(15), A(14) => A1(14), A(13) => 
                           A1(13), A(12) => A1(12), A(11) => A1(11), A(10) => 
                           A1(10), A(9) => A1(9), A(8) => A1(8), A(7) => A1(7),
                           A(6) => A1(6), A(5) => A1(5), A(4) => A1(4), A(3) =>
                           A1(3), A(2) => A1(2), A(1) => A1(1), A(0) => A1(0), 
                           B(15) => A2(15), B(14) => A2(14), B(13) => A2(13), 
                           B(12) => A2(12), B(11) => A2(11), B(10) => A2(10), 
                           B(9) => A2(9), B(8) => A2(8), B(7) => A2(7), B(6) =>
                           A2(6), B(5) => A2(5), B(4) => A2(4), B(3) => A2(3), 
                           B(2) => A2(2), B(1) => A2(1), B(0) => A2(0), S => 
                           S(0), Y(15) => out1_15_port, Y(14) => out1_14_port, 
                           Y(13) => out1_13_port, Y(12) => out1_12_port, Y(11) 
                           => out1_11_port, Y(10) => out1_10_port, Y(9) => 
                           out1_9_port, Y(8) => out1_8_port, Y(7) => 
                           out1_7_port, Y(6) => out1_6_port, Y(5) => 
                           out1_5_port, Y(4) => out1_4_port, Y(3) => 
                           out1_3_port, Y(2) => out1_2_port, Y(1) => 
                           out1_1_port, Y(0) => out1_0_port);
   MUX2 : muxN1_N16_27 port map( A(15) => A3(15), A(14) => A3(14), A(13) => 
                           A3(13), A(12) => A3(12), A(11) => A3(11), A(10) => 
                           A3(10), A(9) => A3(9), A(8) => A3(8), A(7) => A3(7),
                           A(6) => A3(6), A(5) => A3(5), A(4) => A3(4), A(3) =>
                           A3(3), A(2) => A3(2), A(1) => A3(1), A(0) => A3(0), 
                           B(15) => A4(15), B(14) => A4(14), B(13) => A4(13), 
                           B(12) => A4(12), B(11) => A4(11), B(10) => A4(10), 
                           B(9) => A4(9), B(8) => A4(8), B(7) => A4(7), B(6) =>
                           A4(6), B(5) => A4(5), B(4) => A4(4), B(3) => A4(3), 
                           B(2) => A4(2), B(1) => A4(1), B(0) => A4(0), S => 
                           S(0), Y(15) => out2_15_port, Y(14) => out2_14_port, 
                           Y(13) => out2_13_port, Y(12) => out2_12_port, Y(11) 
                           => out2_11_port, Y(10) => out2_10_port, Y(9) => 
                           out2_9_port, Y(8) => out2_8_port, Y(7) => 
                           out2_7_port, Y(6) => out2_6_port, Y(5) => 
                           out2_5_port, Y(4) => out2_4_port, Y(3) => 
                           out2_3_port, Y(2) => out2_2_port, Y(1) => 
                           out2_1_port, Y(0) => out2_0_port);
   MUX3 : muxN1_N16_26 port map( A(15) => A5(15), A(14) => A5(14), A(13) => 
                           A5(13), A(12) => A5(12), A(11) => A5(11), A(10) => 
                           A5(10), A(9) => A5(9), A(8) => A5(8), A(7) => A5(7),
                           A(6) => A5(6), A(5) => A5(5), A(4) => A5(4), A(3) =>
                           A5(3), A(2) => A5(2), A(1) => A5(1), A(0) => A5(0), 
                           B(15) => A6(15), B(14) => A6(14), B(13) => A6(13), 
                           B(12) => A6(12), B(11) => A6(11), B(10) => A6(10), 
                           B(9) => A6(9), B(8) => A6(8), B(7) => A6(7), B(6) =>
                           A6(6), B(5) => A6(5), B(4) => A6(4), B(3) => A6(3), 
                           B(2) => A6(2), B(1) => A6(1), B(0) => A6(0), S => 
                           S(0), Y(15) => out3_15_port, Y(14) => out3_14_port, 
                           Y(13) => out3_13_port, Y(12) => out3_12_port, Y(11) 
                           => out3_11_port, Y(10) => out3_10_port, Y(9) => 
                           out3_9_port, Y(8) => out3_8_port, Y(7) => 
                           out3_7_port, Y(6) => out3_6_port, Y(5) => 
                           out3_5_port, Y(4) => out3_4_port, Y(3) => 
                           out3_3_port, Y(2) => out3_2_port, Y(1) => 
                           out3_1_port, Y(0) => out3_0_port);
   MUX4 : muxN1_N16_25 port map( A(15) => A7(15), A(14) => A7(14), A(13) => 
                           A7(13), A(12) => A7(12), A(11) => A7(11), A(10) => 
                           A7(10), A(9) => A7(9), A(8) => A7(8), A(7) => A7(7),
                           A(6) => A7(6), A(5) => A7(5), A(4) => A7(4), A(3) =>
                           A7(3), A(2) => A7(2), A(1) => A7(1), A(0) => A7(0), 
                           B(15) => A8(15), B(14) => A8(14), B(13) => A8(13), 
                           B(12) => A8(12), B(11) => A8(11), B(10) => A8(10), 
                           B(9) => A8(9), B(8) => A8(8), B(7) => A8(7), B(6) =>
                           A8(6), B(5) => A8(5), B(4) => A8(4), B(3) => A8(3), 
                           B(2) => A8(2), B(1) => A8(1), B(0) => A8(0), S => 
                           S(0), Y(15) => out4_15_port, Y(14) => out4_14_port, 
                           Y(13) => out4_13_port, Y(12) => out4_12_port, Y(11) 
                           => out4_11_port, Y(10) => out4_10_port, Y(9) => 
                           out4_9_port, Y(8) => out4_8_port, Y(7) => 
                           out4_7_port, Y(6) => out4_6_port, Y(5) => 
                           out4_5_port, Y(4) => out4_4_port, Y(3) => 
                           out4_3_port, Y(2) => out4_2_port, Y(1) => 
                           out4_1_port, Y(0) => out4_0_port);
   MUX5 : muxN1_N16_24 port map( A(15) => out1_15_port, A(14) => out1_14_port, 
                           A(13) => out1_13_port, A(12) => out1_12_port, A(11) 
                           => out1_11_port, A(10) => out1_10_port, A(9) => 
                           out1_9_port, A(8) => out1_8_port, A(7) => 
                           out1_7_port, A(6) => out1_6_port, A(5) => 
                           out1_5_port, A(4) => out1_4_port, A(3) => 
                           out1_3_port, A(2) => out1_2_port, A(1) => 
                           out1_1_port, A(0) => out1_0_port, B(15) => 
                           out2_15_port, B(14) => out2_14_port, B(13) => 
                           out2_13_port, B(12) => out2_12_port, B(11) => 
                           out2_11_port, B(10) => out2_10_port, B(9) => 
                           out2_9_port, B(8) => out2_8_port, B(7) => 
                           out2_7_port, B(6) => out2_6_port, B(5) => 
                           out2_5_port, B(4) => out2_4_port, B(3) => 
                           out2_3_port, B(2) => out2_2_port, B(1) => 
                           out2_1_port, B(0) => out2_0_port, S => S(1), Y(15) 
                           => out5_15_port, Y(14) => out5_14_port, Y(13) => 
                           out5_13_port, Y(12) => out5_12_port, Y(11) => 
                           out5_11_port, Y(10) => out5_10_port, Y(9) => 
                           out5_9_port, Y(8) => out5_8_port, Y(7) => 
                           out5_7_port, Y(6) => out5_6_port, Y(5) => 
                           out5_5_port, Y(4) => out5_4_port, Y(3) => 
                           out5_3_port, Y(2) => out5_2_port, Y(1) => 
                           out5_1_port, Y(0) => out5_0_port);
   MUX6 : muxN1_N16_23 port map( A(15) => out3_15_port, A(14) => out3_14_port, 
                           A(13) => out3_13_port, A(12) => out3_12_port, A(11) 
                           => out3_11_port, A(10) => out3_10_port, A(9) => 
                           out3_9_port, A(8) => out3_8_port, A(7) => 
                           out3_7_port, A(6) => out3_6_port, A(5) => 
                           out3_5_port, A(4) => out3_4_port, A(3) => 
                           out3_3_port, A(2) => out3_2_port, A(1) => 
                           out3_1_port, A(0) => out3_0_port, B(15) => 
                           out4_15_port, B(14) => out4_14_port, B(13) => 
                           out4_13_port, B(12) => out4_12_port, B(11) => 
                           out4_11_port, B(10) => out4_10_port, B(9) => 
                           out4_9_port, B(8) => out4_8_port, B(7) => 
                           out4_7_port, B(6) => out4_6_port, B(5) => 
                           out4_5_port, B(4) => out4_4_port, B(3) => 
                           out4_3_port, B(2) => out4_2_port, B(1) => 
                           out4_1_port, B(0) => out4_0_port, S => S(1), Y(15) 
                           => out6_15_port, Y(14) => out6_14_port, Y(13) => 
                           out6_13_port, Y(12) => out6_12_port, Y(11) => 
                           out6_11_port, Y(10) => out6_10_port, Y(9) => 
                           out6_9_port, Y(8) => out6_8_port, Y(7) => 
                           out6_7_port, Y(6) => out6_6_port, Y(5) => 
                           out6_5_port, Y(4) => out6_4_port, Y(3) => 
                           out6_3_port, Y(2) => out6_2_port, Y(1) => 
                           out6_1_port, Y(0) => out6_0_port);
   MUX7 : muxN1_N16_22 port map( A(15) => out5_15_port, A(14) => out5_14_port, 
                           A(13) => out5_13_port, A(12) => out5_12_port, A(11) 
                           => out5_11_port, A(10) => out5_10_port, A(9) => 
                           out5_9_port, A(8) => out5_8_port, A(7) => 
                           out5_7_port, A(6) => out5_6_port, A(5) => 
                           out5_5_port, A(4) => out5_4_port, A(3) => 
                           out5_3_port, A(2) => out5_2_port, A(1) => 
                           out5_1_port, A(0) => out5_0_port, B(15) => 
                           out6_15_port, B(14) => out6_14_port, B(13) => 
                           out6_13_port, B(12) => out6_12_port, B(11) => 
                           out6_11_port, B(10) => out6_10_port, B(9) => 
                           out6_9_port, B(8) => out6_8_port, B(7) => 
                           out6_7_port, B(6) => out6_6_port, B(5) => 
                           out6_5_port, B(4) => out6_4_port, B(3) => 
                           out6_3_port, B(2) => out6_2_port, B(1) => 
                           out6_1_port, B(0) => out6_0_port, S => S(2), Y(15) 
                           => Y(15), Y(14) => Y(14), Y(13) => Y(13), Y(12) => 
                           Y(12), Y(11) => Y(11), Y(10) => Y(10), Y(9) => Y(9),
                           Y(8) => Y(8), Y(7) => Y(7), Y(6) => Y(6), Y(5) => 
                           Y(5), Y(4) => Y(4), Y(3) => Y(3), Y(2) => Y(2), Y(1)
                           => Y(1), Y(0) => Y(0));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity complementor_N16_0 is

   port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (15 
         downto 0));

end complementor_N16_0;

architecture SYN_ARCHDATAFLOW of complementor_N16_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component complementor_N16_0_DW01_inc_0_DW01_inc_7
      port( A : in std_logic_vector (15 downto 0);  SUM : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal N9, N8, N7, N6, N5, N4, N3, N2, N15, N14, N13, N12, N11, N10, N1, N0 
      : std_logic;

begin
   
   add_0_root_add_19_ni : complementor_N16_0_DW01_inc_0_DW01_inc_7 port map( 
                           A(15) => N0, A(14) => N1, A(13) => N2, A(12) => N3, 
                           A(11) => N4, A(10) => N5, A(9) => N6, A(8) => N7, 
                           A(7) => N8, A(6) => N9, A(5) => N10, A(4) => N11, 
                           A(3) => N12, A(2) => N13, A(1) => N14, A(0) => N15, 
                           SUM(15) => Y(15), SUM(14) => Y(14), SUM(13) => Y(13)
                           , SUM(12) => Y(12), SUM(11) => Y(11), SUM(10) => 
                           Y(10), SUM(9) => Y(9), SUM(8) => Y(8), SUM(7) => 
                           Y(7), SUM(6) => Y(6), SUM(5) => Y(5), SUM(4) => Y(4)
                           , SUM(3) => Y(3), SUM(2) => Y(2), SUM(1) => Y(1), 
                           SUM(0) => Y(0));
   U2 : INV_X1 port map( A => A(6), ZN => N9);
   U3 : INV_X1 port map( A => A(7), ZN => N8);
   U4 : INV_X1 port map( A => A(8), ZN => N7);
   U5 : INV_X1 port map( A => A(9), ZN => N6);
   U6 : INV_X1 port map( A => A(10), ZN => N5);
   U7 : INV_X1 port map( A => A(11), ZN => N4);
   U8 : INV_X1 port map( A => A(12), ZN => N3);
   U9 : INV_X1 port map( A => A(13), ZN => N2);
   U10 : INV_X1 port map( A => A(0), ZN => N15);
   U11 : INV_X1 port map( A => A(1), ZN => N14);
   U12 : INV_X1 port map( A => A(2), ZN => N13);
   U13 : INV_X1 port map( A => A(3), ZN => N12);
   U14 : INV_X1 port map( A => A(4), ZN => N11);
   U15 : INV_X1 port map( A => A(5), ZN => N10);
   U16 : INV_X1 port map( A => A(14), ZN => N1);
   U17 : INV_X1 port map( A => A(15), ZN => N0);

end SYN_ARCHDATAFLOW;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity shift_pow2_N8_0 is

   port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector (3 
         downto 0);  SA : out std_logic_vector (15 downto 0));

end shift_pow2_N8_0;

architecture SYN_ARCHBEH of shift_pow2_N8_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component shift_pow2_N8_0_DW02_mult_0_DW02_mult_7
      port( A, B : in std_logic_vector (7 downto 0);  TC : in std_logic;  
            PRODUCT : out std_logic_vector (15 downto 0));
   end component;
   
   signal n4, shift_pow_31_ML_int_4_0_port, shift_pow_31_ML_int_4_1_port, 
      shift_pow_31_ML_int_4_2_port, shift_pow_31_ML_int_4_3_port, 
      shift_pow_31_ML_int_4_4_port, shift_pow_31_ML_int_4_5_port, 
      shift_pow_31_ML_int_4_6_port, shift_pow_31_ML_int_4_7_port, 
      shift_pow_31_ML_int_2_0_port, shift_pow_31_ML_int_2_1_port, n1, n2, n3, 
      n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   n4 <= '0';
   mult_31 : shift_pow2_N8_0_DW02_mult_0_DW02_mult_7 port map( A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), B(7)
                           => shift_pow_31_ML_int_4_7_port, B(6) => 
                           shift_pow_31_ML_int_4_6_port, B(5) => 
                           shift_pow_31_ML_int_4_5_port, B(4) => 
                           shift_pow_31_ML_int_4_4_port, B(3) => 
                           shift_pow_31_ML_int_4_3_port, B(2) => 
                           shift_pow_31_ML_int_4_2_port, B(1) => 
                           shift_pow_31_ML_int_4_1_port, B(0) => 
                           shift_pow_31_ML_int_4_0_port, TC => n4, PRODUCT(15) 
                           => SA(15), PRODUCT(14) => SA(14), PRODUCT(13) => 
                           SA(13), PRODUCT(12) => SA(12), PRODUCT(11) => SA(11)
                           , PRODUCT(10) => SA(10), PRODUCT(9) => SA(9), 
                           PRODUCT(8) => SA(8), PRODUCT(7) => SA(7), PRODUCT(6)
                           => SA(6), PRODUCT(5) => SA(5), PRODUCT(4) => SA(4), 
                           PRODUCT(3) => SA(3), PRODUCT(2) => SA(2), PRODUCT(1)
                           => SA(1), PRODUCT(0) => SA(0));
   U3 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_1_port, 
                           ZN => n1);
   U4 : AND2_X1 port map( A1 => Shift(2), A2 => shift_pow_31_ML_int_2_0_port, 
                           ZN => n2);
   U5 : AND2_X1 port map( A1 => Shift(2), A2 => n6, ZN => n3);
   U7 : AND2_X1 port map( A1 => Shift(2), A2 => n7, ZN => n5);
   U8 : AND2_X1 port map( A1 => Shift(1), A2 => n10, ZN => n6);
   U9 : AND2_X1 port map( A1 => Shift(1), A2 => Shift(0), ZN => n7);
   U10 : AND2_X1 port map( A1 => n5, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_7_port);
   U11 : AND2_X1 port map( A1 => n3, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_6_port);
   U12 : AND2_X1 port map( A1 => n1, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_5_port);
   U13 : AND2_X1 port map( A1 => n2, A2 => n8, ZN => 
                           shift_pow_31_ML_int_4_4_port);
   U14 : INV_X1 port map( A => Shift(3), ZN => n8);
   U15 : AND2_X1 port map( A1 => n7, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_3_port);
   U16 : AND2_X1 port map( A1 => n6, A2 => n9, ZN => 
                           shift_pow_31_ML_int_4_2_port);
   U17 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_1_port, ZN => 
                           shift_pow_31_ML_int_4_1_port);
   U18 : AND2_X1 port map( A1 => n9, A2 => shift_pow_31_ML_int_2_0_port, ZN => 
                           shift_pow_31_ML_int_4_0_port);
   U19 : NOR2_X1 port map( A1 => Shift(3), A2 => Shift(2), ZN => n9);
   U20 : NOR2_X1 port map( A1 => n10, A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_1_port);
   U21 : NOR2_X1 port map( A1 => Shift(0), A2 => Shift(1), ZN => 
                           shift_pow_31_ML_int_2_0_port);
   U22 : INV_X1 port map( A => Shift(0), ZN => n10);

end SYN_ARCHBEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity booth_encoder_N8 is

   port( B : in std_logic_vector (7 downto 0);  S : out std_logic_vector (11 
         downto 0));

end booth_encoder_N8;

architecture SYN_ARCHSTRUCT of booth_encoder_N8 is

   component booth_encoder_block_17
      port( Bi : in std_logic_vector (2 downto 0);  So : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component booth_encoder_block_18
      port( Bi : in std_logic_vector (2 downto 0);  So : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component booth_encoder_block_19
      port( Bi : in std_logic_vector (2 downto 0);  So : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component booth_encoder_block_16
      port( Bi : in std_logic_vector (2 downto 0);  So : out std_logic_vector 
            (2 downto 0));
   end component;
   
   signal X_Logic0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   BLK_0 : booth_encoder_block_16 port map( Bi(2) => B(1), Bi(1) => B(0), Bi(0)
                           => X_Logic0_port, So(2) => S(2), So(1) => S(1), 
                           So(0) => S(0));
   BLK_1 : booth_encoder_block_19 port map( Bi(2) => B(3), Bi(1) => B(2), Bi(0)
                           => B(1), So(2) => S(5), So(1) => S(4), So(0) => S(3)
                           );
   BLK_2 : booth_encoder_block_18 port map( Bi(2) => B(5), Bi(1) => B(4), Bi(0)
                           => B(3), So(2) => S(8), So(1) => S(7), So(0) => S(6)
                           );
   BLK_3 : booth_encoder_block_17 port map( Bi(2) => B(7), Bi(1) => B(6), Bi(0)
                           => B(5), So(2) => S(11), So(1) => S(10), So(0) => 
                           S(9));

end SYN_ARCHSTRUCT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N8.all;

entity BOOTHMUL_N8 is

   port( A, B : in std_logic_vector (7 downto 0);  Y : out std_logic_vector (15
         downto 0));

end BOOTHMUL_N8;

architecture SYN_ARCHSTRUCT of BOOTHMUL_N8 is

   component P4_adder_N16_Nbit_blocks4_1
      port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (15 downto 0);  Cout : out std_logic);
   end component;
   
   component P4_adder_N16_Nbit_blocks4_2
      port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (15 downto 0);  Cout : out std_logic);
   end component;
   
   component P4_adder_N16_Nbit_blocks4_0
      port( A, B : in std_logic_vector (15 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (15 downto 0);  Cout : out std_logic);
   end component;
   
   component mux_8to1_N16_1
      port( A1, A2, A3, A4, A5, A6, A7, A8 : in std_logic_vector (15 downto 0);
            S : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (15
            downto 0));
   end component;
   
   component mux_8to1_N16_2
      port( A1, A2, A3, A4, A5, A6, A7, A8 : in std_logic_vector (15 downto 0);
            S : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (15
            downto 0));
   end component;
   
   component mux_8to1_N16_3
      port( A1, A2, A3, A4, A5, A6, A7, A8 : in std_logic_vector (15 downto 0);
            S : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (15
            downto 0));
   end component;
   
   component mux_8to1_N16_0
      port( A1, A2, A3, A4, A5, A6, A7, A8 : in std_logic_vector (15 downto 0);
            S : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (15
            downto 0));
   end component;
   
   component complementor_N16_1
      port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component complementor_N16_2
      port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component complementor_N16_3
      port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component complementor_N16_4
      port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component complementor_N16_5
      port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component complementor_N16_6
      port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component complementor_N16_7
      port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component complementor_N16_0
      port( A : in std_logic_vector (15 downto 0);  Y : out std_logic_vector 
            (15 downto 0));
   end component;
   
   component shift_pow2_N8_1
      port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector 
            (3 downto 0);  SA : out std_logic_vector (15 downto 0));
   end component;
   
   component shift_pow2_N8_2
      port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector 
            (3 downto 0);  SA : out std_logic_vector (15 downto 0));
   end component;
   
   component shift_pow2_N8_3
      port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector 
            (3 downto 0);  SA : out std_logic_vector (15 downto 0));
   end component;
   
   component shift_pow2_N8_4
      port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector 
            (3 downto 0);  SA : out std_logic_vector (15 downto 0));
   end component;
   
   component shift_pow2_N8_5
      port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector 
            (3 downto 0);  SA : out std_logic_vector (15 downto 0));
   end component;
   
   component shift_pow2_N8_6
      port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector 
            (3 downto 0);  SA : out std_logic_vector (15 downto 0));
   end component;
   
   component shift_pow2_N8_7
      port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector 
            (3 downto 0);  SA : out std_logic_vector (15 downto 0));
   end component;
   
   component shift_pow2_N8_0
      port( A : in std_logic_vector (7 downto 0);  Shift : in std_logic_vector 
            (3 downto 0);  SA : out std_logic_vector (15 downto 0));
   end component;
   
   component booth_encoder_N8
      port( B : in std_logic_vector (7 downto 0);  S : out std_logic_vector (11
            downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sel_muxes_11_port, sel_muxes_10_port, 
      sel_muxes_9_port, sel_muxes_8_port, sel_muxes_7_port, sel_muxes_6_port, 
      sel_muxes_5_port, sel_muxes_4_port, sel_muxes_3_port, sel_muxes_2_port, 
      sel_muxes_1_port, sel_muxes_0_port, out_shifter_7_15_port, 
      out_shifter_7_14_port, out_shifter_7_13_port, out_shifter_7_12_port, 
      out_shifter_7_11_port, out_shifter_7_10_port, out_shifter_7_9_port, 
      out_shifter_7_8_port, out_shifter_7_7_port, out_shifter_7_6_port, 
      out_shifter_7_5_port, out_shifter_7_4_port, out_shifter_7_3_port, 
      out_shifter_7_2_port, out_shifter_7_1_port, out_shifter_7_0_port, 
      out_shifter_6_15_port, out_shifter_6_14_port, out_shifter_6_13_port, 
      out_shifter_6_12_port, out_shifter_6_11_port, out_shifter_6_10_port, 
      out_shifter_6_9_port, out_shifter_6_8_port, out_shifter_6_7_port, 
      out_shifter_6_6_port, out_shifter_6_5_port, out_shifter_6_4_port, 
      out_shifter_6_3_port, out_shifter_6_2_port, out_shifter_6_1_port, 
      out_shifter_6_0_port, out_shifter_5_15_port, out_shifter_5_14_port, 
      out_shifter_5_13_port, out_shifter_5_12_port, out_shifter_5_11_port, 
      out_shifter_5_10_port, out_shifter_5_9_port, out_shifter_5_8_port, 
      out_shifter_5_7_port, out_shifter_5_6_port, out_shifter_5_5_port, 
      out_shifter_5_4_port, out_shifter_5_3_port, out_shifter_5_2_port, 
      out_shifter_5_1_port, out_shifter_5_0_port, out_shifter_4_15_port, 
      out_shifter_4_14_port, out_shifter_4_13_port, out_shifter_4_12_port, 
      out_shifter_4_11_port, out_shifter_4_10_port, out_shifter_4_9_port, 
      out_shifter_4_8_port, out_shifter_4_7_port, out_shifter_4_6_port, 
      out_shifter_4_5_port, out_shifter_4_4_port, out_shifter_4_3_port, 
      out_shifter_4_2_port, out_shifter_4_1_port, out_shifter_4_0_port, 
      out_shifter_3_15_port, out_shifter_3_14_port, out_shifter_3_13_port, 
      out_shifter_3_12_port, out_shifter_3_11_port, out_shifter_3_10_port, 
      out_shifter_3_9_port, out_shifter_3_8_port, out_shifter_3_7_port, 
      out_shifter_3_6_port, out_shifter_3_5_port, out_shifter_3_4_port, 
      out_shifter_3_3_port, out_shifter_3_2_port, out_shifter_3_1_port, 
      out_shifter_3_0_port, out_shifter_2_15_port, out_shifter_2_14_port, 
      out_shifter_2_13_port, out_shifter_2_12_port, out_shifter_2_11_port, 
      out_shifter_2_10_port, out_shifter_2_9_port, out_shifter_2_8_port, 
      out_shifter_2_7_port, out_shifter_2_6_port, out_shifter_2_5_port, 
      out_shifter_2_4_port, out_shifter_2_3_port, out_shifter_2_2_port, 
      out_shifter_2_1_port, out_shifter_2_0_port, out_shifter_1_15_port, 
      out_shifter_1_14_port, out_shifter_1_13_port, out_shifter_1_12_port, 
      out_shifter_1_11_port, out_shifter_1_10_port, out_shifter_1_9_port, 
      out_shifter_1_8_port, out_shifter_1_7_port, out_shifter_1_6_port, 
      out_shifter_1_5_port, out_shifter_1_4_port, out_shifter_1_3_port, 
      out_shifter_1_2_port, out_shifter_1_1_port, out_shifter_1_0_port, 
      out_shifter_0_15_port, out_shifter_0_14_port, out_shifter_0_13_port, 
      out_shifter_0_12_port, out_shifter_0_11_port, out_shifter_0_10_port, 
      out_shifter_0_9_port, out_shifter_0_8_port, out_shifter_0_7_port, 
      out_shifter_0_6_port, out_shifter_0_5_port, out_shifter_0_4_port, 
      out_shifter_0_3_port, out_shifter_0_2_port, out_shifter_0_1_port, 
      out_shifter_0_0_port, out_shifter_neg_7_15_port, 
      out_shifter_neg_7_14_port, out_shifter_neg_7_13_port, 
      out_shifter_neg_7_12_port, out_shifter_neg_7_11_port, 
      out_shifter_neg_7_10_port, out_shifter_neg_7_9_port, 
      out_shifter_neg_7_8_port, out_shifter_neg_7_7_port, 
      out_shifter_neg_7_6_port, out_shifter_neg_7_5_port, 
      out_shifter_neg_7_4_port, out_shifter_neg_7_3_port, 
      out_shifter_neg_7_2_port, out_shifter_neg_7_1_port, 
      out_shifter_neg_7_0_port, out_shifter_neg_6_15_port, 
      out_shifter_neg_6_14_port, out_shifter_neg_6_13_port, 
      out_shifter_neg_6_12_port, out_shifter_neg_6_11_port, 
      out_shifter_neg_6_10_port, out_shifter_neg_6_9_port, 
      out_shifter_neg_6_8_port, out_shifter_neg_6_7_port, 
      out_shifter_neg_6_6_port, out_shifter_neg_6_5_port, 
      out_shifter_neg_6_4_port, out_shifter_neg_6_3_port, 
      out_shifter_neg_6_2_port, out_shifter_neg_6_1_port, 
      out_shifter_neg_6_0_port, out_shifter_neg_5_15_port, 
      out_shifter_neg_5_14_port, out_shifter_neg_5_13_port, 
      out_shifter_neg_5_12_port, out_shifter_neg_5_11_port, 
      out_shifter_neg_5_10_port, out_shifter_neg_5_9_port, 
      out_shifter_neg_5_8_port, out_shifter_neg_5_7_port, 
      out_shifter_neg_5_6_port, out_shifter_neg_5_5_port, 
      out_shifter_neg_5_4_port, out_shifter_neg_5_3_port, 
      out_shifter_neg_5_2_port, out_shifter_neg_5_1_port, 
      out_shifter_neg_5_0_port, out_shifter_neg_4_15_port, 
      out_shifter_neg_4_14_port, out_shifter_neg_4_13_port, 
      out_shifter_neg_4_12_port, out_shifter_neg_4_11_port, 
      out_shifter_neg_4_10_port, out_shifter_neg_4_9_port, 
      out_shifter_neg_4_8_port, out_shifter_neg_4_7_port, 
      out_shifter_neg_4_6_port, out_shifter_neg_4_5_port, 
      out_shifter_neg_4_4_port, out_shifter_neg_4_3_port, 
      out_shifter_neg_4_2_port, out_shifter_neg_4_1_port, 
      out_shifter_neg_4_0_port, out_shifter_neg_3_15_port, 
      out_shifter_neg_3_14_port, out_shifter_neg_3_13_port, 
      out_shifter_neg_3_12_port, out_shifter_neg_3_11_port, 
      out_shifter_neg_3_10_port, out_shifter_neg_3_9_port, 
      out_shifter_neg_3_8_port, out_shifter_neg_3_7_port, 
      out_shifter_neg_3_6_port, out_shifter_neg_3_5_port, 
      out_shifter_neg_3_4_port, out_shifter_neg_3_3_port, 
      out_shifter_neg_3_2_port, out_shifter_neg_3_1_port, 
      out_shifter_neg_3_0_port, out_shifter_neg_2_15_port, 
      out_shifter_neg_2_14_port, out_shifter_neg_2_13_port, 
      out_shifter_neg_2_12_port, out_shifter_neg_2_11_port, 
      out_shifter_neg_2_10_port, out_shifter_neg_2_9_port, 
      out_shifter_neg_2_8_port, out_shifter_neg_2_7_port, 
      out_shifter_neg_2_6_port, out_shifter_neg_2_5_port, 
      out_shifter_neg_2_4_port, out_shifter_neg_2_3_port, 
      out_shifter_neg_2_2_port, out_shifter_neg_2_1_port, 
      out_shifter_neg_2_0_port, out_shifter_neg_1_15_port, 
      out_shifter_neg_1_14_port, out_shifter_neg_1_13_port, 
      out_shifter_neg_1_12_port, out_shifter_neg_1_11_port, 
      out_shifter_neg_1_10_port, out_shifter_neg_1_9_port, 
      out_shifter_neg_1_8_port, out_shifter_neg_1_7_port, 
      out_shifter_neg_1_6_port, out_shifter_neg_1_5_port, 
      out_shifter_neg_1_4_port, out_shifter_neg_1_3_port, 
      out_shifter_neg_1_2_port, out_shifter_neg_1_1_port, 
      out_shifter_neg_1_0_port, out_shifter_neg_0_15_port, 
      out_shifter_neg_0_14_port, out_shifter_neg_0_13_port, 
      out_shifter_neg_0_12_port, out_shifter_neg_0_11_port, 
      out_shifter_neg_0_10_port, out_shifter_neg_0_9_port, 
      out_shifter_neg_0_8_port, out_shifter_neg_0_7_port, 
      out_shifter_neg_0_6_port, out_shifter_neg_0_5_port, 
      out_shifter_neg_0_4_port, out_shifter_neg_0_3_port, 
      out_shifter_neg_0_2_port, out_shifter_neg_0_1_port, 
      out_shifter_neg_0_0_port, out_muxes_3_15_port, out_muxes_3_14_port, 
      out_muxes_3_13_port, out_muxes_3_12_port, out_muxes_3_11_port, 
      out_muxes_3_10_port, out_muxes_3_9_port, out_muxes_3_8_port, 
      out_muxes_3_7_port, out_muxes_3_6_port, out_muxes_3_5_port, 
      out_muxes_3_4_port, out_muxes_3_3_port, out_muxes_3_2_port, 
      out_muxes_3_1_port, out_muxes_3_0_port, out_muxes_2_15_port, 
      out_muxes_2_14_port, out_muxes_2_13_port, out_muxes_2_12_port, 
      out_muxes_2_11_port, out_muxes_2_10_port, out_muxes_2_9_port, 
      out_muxes_2_8_port, out_muxes_2_7_port, out_muxes_2_6_port, 
      out_muxes_2_5_port, out_muxes_2_4_port, out_muxes_2_3_port, 
      out_muxes_2_2_port, out_muxes_2_1_port, out_muxes_2_0_port, 
      out_muxes_1_15_port, out_muxes_1_14_port, out_muxes_1_13_port, 
      out_muxes_1_12_port, out_muxes_1_11_port, out_muxes_1_10_port, 
      out_muxes_1_9_port, out_muxes_1_8_port, out_muxes_1_7_port, 
      out_muxes_1_6_port, out_muxes_1_5_port, out_muxes_1_4_port, 
      out_muxes_1_3_port, out_muxes_1_2_port, out_muxes_1_1_port, 
      out_muxes_1_0_port, out_muxes_0_15_port, out_muxes_0_14_port, 
      out_muxes_0_13_port, out_muxes_0_12_port, out_muxes_0_11_port, 
      out_muxes_0_10_port, out_muxes_0_9_port, out_muxes_0_8_port, 
      out_muxes_0_7_port, out_muxes_0_6_port, out_muxes_0_5_port, 
      out_muxes_0_4_port, out_muxes_0_3_port, out_muxes_0_2_port, 
      out_muxes_0_1_port, out_muxes_0_0_port, out_adder_1_15_port, 
      out_adder_1_14_port, out_adder_1_13_port, out_adder_1_12_port, 
      out_adder_1_11_port, out_adder_1_10_port, out_adder_1_9_port, 
      out_adder_1_8_port, out_adder_1_7_port, out_adder_1_6_port, 
      out_adder_1_5_port, out_adder_1_4_port, out_adder_1_3_port, 
      out_adder_1_2_port, out_adder_1_1_port, out_adder_1_0_port, 
      out_adder_0_15_port, out_adder_0_14_port, out_adder_0_13_port, 
      out_adder_0_12_port, out_adder_0_11_port, out_adder_0_10_port, 
      out_adder_0_9_port, out_adder_0_8_port, out_adder_0_7_port, 
      out_adder_0_6_port, out_adder_0_5_port, out_adder_0_4_port, 
      out_adder_0_3_port, out_adder_0_2_port, out_adder_0_1_port, 
      out_adder_0_0_port, n_1123, n_1124, n_1125 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   BE : booth_encoder_N8 port map( B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), S(11) => sel_muxes_11_port, 
                           S(10) => sel_muxes_10_port, S(9) => sel_muxes_9_port
                           , S(8) => sel_muxes_8_port, S(7) => sel_muxes_7_port
                           , S(6) => sel_muxes_6_port, S(5) => sel_muxes_5_port
                           , S(4) => sel_muxes_4_port, S(3) => sel_muxes_3_port
                           , S(2) => sel_muxes_2_port, S(1) => sel_muxes_1_port
                           , S(0) => sel_muxes_0_port);
   SHFT_0 : shift_pow2_N8_0 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5),
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), Shift(3) => X_Logic0_port, 
                           Shift(2) => X_Logic0_port, Shift(1) => X_Logic0_port
                           , Shift(0) => X_Logic0_port, SA(15) => 
                           out_shifter_0_15_port, SA(14) => 
                           out_shifter_0_14_port, SA(13) => 
                           out_shifter_0_13_port, SA(12) => 
                           out_shifter_0_12_port, SA(11) => 
                           out_shifter_0_11_port, SA(10) => 
                           out_shifter_0_10_port, SA(9) => out_shifter_0_9_port
                           , SA(8) => out_shifter_0_8_port, SA(7) => 
                           out_shifter_0_7_port, SA(6) => out_shifter_0_6_port,
                           SA(5) => out_shifter_0_5_port, SA(4) => 
                           out_shifter_0_4_port, SA(3) => out_shifter_0_3_port,
                           SA(2) => out_shifter_0_2_port, SA(1) => 
                           out_shifter_0_1_port, SA(0) => out_shifter_0_0_port)
                           ;
   SHFT_1 : shift_pow2_N8_7 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5),
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), Shift(3) => X_Logic0_port, 
                           Shift(2) => X_Logic0_port, Shift(1) => X_Logic0_port
                           , Shift(0) => X_Logic1_port, SA(15) => 
                           out_shifter_1_15_port, SA(14) => 
                           out_shifter_1_14_port, SA(13) => 
                           out_shifter_1_13_port, SA(12) => 
                           out_shifter_1_12_port, SA(11) => 
                           out_shifter_1_11_port, SA(10) => 
                           out_shifter_1_10_port, SA(9) => out_shifter_1_9_port
                           , SA(8) => out_shifter_1_8_port, SA(7) => 
                           out_shifter_1_7_port, SA(6) => out_shifter_1_6_port,
                           SA(5) => out_shifter_1_5_port, SA(4) => 
                           out_shifter_1_4_port, SA(3) => out_shifter_1_3_port,
                           SA(2) => out_shifter_1_2_port, SA(1) => 
                           out_shifter_1_1_port, SA(0) => out_shifter_1_0_port)
                           ;
   SHFT_2 : shift_pow2_N8_6 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5),
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), Shift(3) => X_Logic0_port, 
                           Shift(2) => X_Logic0_port, Shift(1) => X_Logic1_port
                           , Shift(0) => X_Logic0_port, SA(15) => 
                           out_shifter_2_15_port, SA(14) => 
                           out_shifter_2_14_port, SA(13) => 
                           out_shifter_2_13_port, SA(12) => 
                           out_shifter_2_12_port, SA(11) => 
                           out_shifter_2_11_port, SA(10) => 
                           out_shifter_2_10_port, SA(9) => out_shifter_2_9_port
                           , SA(8) => out_shifter_2_8_port, SA(7) => 
                           out_shifter_2_7_port, SA(6) => out_shifter_2_6_port,
                           SA(5) => out_shifter_2_5_port, SA(4) => 
                           out_shifter_2_4_port, SA(3) => out_shifter_2_3_port,
                           SA(2) => out_shifter_2_2_port, SA(1) => 
                           out_shifter_2_1_port, SA(0) => out_shifter_2_0_port)
                           ;
   SHFT_3 : shift_pow2_N8_5 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5),
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), Shift(3) => X_Logic0_port, 
                           Shift(2) => X_Logic0_port, Shift(1) => X_Logic1_port
                           , Shift(0) => X_Logic1_port, SA(15) => 
                           out_shifter_3_15_port, SA(14) => 
                           out_shifter_3_14_port, SA(13) => 
                           out_shifter_3_13_port, SA(12) => 
                           out_shifter_3_12_port, SA(11) => 
                           out_shifter_3_11_port, SA(10) => 
                           out_shifter_3_10_port, SA(9) => out_shifter_3_9_port
                           , SA(8) => out_shifter_3_8_port, SA(7) => 
                           out_shifter_3_7_port, SA(6) => out_shifter_3_6_port,
                           SA(5) => out_shifter_3_5_port, SA(4) => 
                           out_shifter_3_4_port, SA(3) => out_shifter_3_3_port,
                           SA(2) => out_shifter_3_2_port, SA(1) => 
                           out_shifter_3_1_port, SA(0) => out_shifter_3_0_port)
                           ;
   SHFT_4 : shift_pow2_N8_4 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5),
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), Shift(3) => X_Logic0_port, 
                           Shift(2) => X_Logic1_port, Shift(1) => X_Logic0_port
                           , Shift(0) => X_Logic0_port, SA(15) => 
                           out_shifter_4_15_port, SA(14) => 
                           out_shifter_4_14_port, SA(13) => 
                           out_shifter_4_13_port, SA(12) => 
                           out_shifter_4_12_port, SA(11) => 
                           out_shifter_4_11_port, SA(10) => 
                           out_shifter_4_10_port, SA(9) => out_shifter_4_9_port
                           , SA(8) => out_shifter_4_8_port, SA(7) => 
                           out_shifter_4_7_port, SA(6) => out_shifter_4_6_port,
                           SA(5) => out_shifter_4_5_port, SA(4) => 
                           out_shifter_4_4_port, SA(3) => out_shifter_4_3_port,
                           SA(2) => out_shifter_4_2_port, SA(1) => 
                           out_shifter_4_1_port, SA(0) => out_shifter_4_0_port)
                           ;
   SHFT_5 : shift_pow2_N8_3 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5),
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), Shift(3) => X_Logic0_port, 
                           Shift(2) => X_Logic1_port, Shift(1) => X_Logic0_port
                           , Shift(0) => X_Logic1_port, SA(15) => 
                           out_shifter_5_15_port, SA(14) => 
                           out_shifter_5_14_port, SA(13) => 
                           out_shifter_5_13_port, SA(12) => 
                           out_shifter_5_12_port, SA(11) => 
                           out_shifter_5_11_port, SA(10) => 
                           out_shifter_5_10_port, SA(9) => out_shifter_5_9_port
                           , SA(8) => out_shifter_5_8_port, SA(7) => 
                           out_shifter_5_7_port, SA(6) => out_shifter_5_6_port,
                           SA(5) => out_shifter_5_5_port, SA(4) => 
                           out_shifter_5_4_port, SA(3) => out_shifter_5_3_port,
                           SA(2) => out_shifter_5_2_port, SA(1) => 
                           out_shifter_5_1_port, SA(0) => out_shifter_5_0_port)
                           ;
   SHFT_6 : shift_pow2_N8_2 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5),
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), Shift(3) => X_Logic0_port, 
                           Shift(2) => X_Logic1_port, Shift(1) => X_Logic1_port
                           , Shift(0) => X_Logic0_port, SA(15) => 
                           out_shifter_6_15_port, SA(14) => 
                           out_shifter_6_14_port, SA(13) => 
                           out_shifter_6_13_port, SA(12) => 
                           out_shifter_6_12_port, SA(11) => 
                           out_shifter_6_11_port, SA(10) => 
                           out_shifter_6_10_port, SA(9) => out_shifter_6_9_port
                           , SA(8) => out_shifter_6_8_port, SA(7) => 
                           out_shifter_6_7_port, SA(6) => out_shifter_6_6_port,
                           SA(5) => out_shifter_6_5_port, SA(4) => 
                           out_shifter_6_4_port, SA(3) => out_shifter_6_3_port,
                           SA(2) => out_shifter_6_2_port, SA(1) => 
                           out_shifter_6_1_port, SA(0) => out_shifter_6_0_port)
                           ;
   SHFT_7 : shift_pow2_N8_1 port map( A(7) => A(7), A(6) => A(6), A(5) => A(5),
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), Shift(3) => X_Logic0_port, 
                           Shift(2) => X_Logic1_port, Shift(1) => X_Logic1_port
                           , Shift(0) => X_Logic1_port, SA(15) => 
                           out_shifter_7_15_port, SA(14) => 
                           out_shifter_7_14_port, SA(13) => 
                           out_shifter_7_13_port, SA(12) => 
                           out_shifter_7_12_port, SA(11) => 
                           out_shifter_7_11_port, SA(10) => 
                           out_shifter_7_10_port, SA(9) => out_shifter_7_9_port
                           , SA(8) => out_shifter_7_8_port, SA(7) => 
                           out_shifter_7_7_port, SA(6) => out_shifter_7_6_port,
                           SA(5) => out_shifter_7_5_port, SA(4) => 
                           out_shifter_7_4_port, SA(3) => out_shifter_7_3_port,
                           SA(2) => out_shifter_7_2_port, SA(1) => 
                           out_shifter_7_1_port, SA(0) => out_shifter_7_0_port)
                           ;
   COMP_0 : complementor_N16_0 port map( A(15) => out_shifter_0_15_port, A(14) 
                           => out_shifter_0_14_port, A(13) => 
                           out_shifter_0_13_port, A(12) => 
                           out_shifter_0_12_port, A(11) => 
                           out_shifter_0_11_port, A(10) => 
                           out_shifter_0_10_port, A(9) => out_shifter_0_9_port,
                           A(8) => out_shifter_0_8_port, A(7) => 
                           out_shifter_0_7_port, A(6) => out_shifter_0_6_port, 
                           A(5) => out_shifter_0_5_port, A(4) => 
                           out_shifter_0_4_port, A(3) => out_shifter_0_3_port, 
                           A(2) => out_shifter_0_2_port, A(1) => 
                           out_shifter_0_1_port, A(0) => out_shifter_0_0_port, 
                           Y(15) => out_shifter_neg_0_15_port, Y(14) => 
                           out_shifter_neg_0_14_port, Y(13) => 
                           out_shifter_neg_0_13_port, Y(12) => 
                           out_shifter_neg_0_12_port, Y(11) => 
                           out_shifter_neg_0_11_port, Y(10) => 
                           out_shifter_neg_0_10_port, Y(9) => 
                           out_shifter_neg_0_9_port, Y(8) => 
                           out_shifter_neg_0_8_port, Y(7) => 
                           out_shifter_neg_0_7_port, Y(6) => 
                           out_shifter_neg_0_6_port, Y(5) => 
                           out_shifter_neg_0_5_port, Y(4) => 
                           out_shifter_neg_0_4_port, Y(3) => 
                           out_shifter_neg_0_3_port, Y(2) => 
                           out_shifter_neg_0_2_port, Y(1) => 
                           out_shifter_neg_0_1_port, Y(0) => 
                           out_shifter_neg_0_0_port);
   COMP_1 : complementor_N16_7 port map( A(15) => out_shifter_1_15_port, A(14) 
                           => out_shifter_1_14_port, A(13) => 
                           out_shifter_1_13_port, A(12) => 
                           out_shifter_1_12_port, A(11) => 
                           out_shifter_1_11_port, A(10) => 
                           out_shifter_1_10_port, A(9) => out_shifter_1_9_port,
                           A(8) => out_shifter_1_8_port, A(7) => 
                           out_shifter_1_7_port, A(6) => out_shifter_1_6_port, 
                           A(5) => out_shifter_1_5_port, A(4) => 
                           out_shifter_1_4_port, A(3) => out_shifter_1_3_port, 
                           A(2) => out_shifter_1_2_port, A(1) => 
                           out_shifter_1_1_port, A(0) => out_shifter_1_0_port, 
                           Y(15) => out_shifter_neg_1_15_port, Y(14) => 
                           out_shifter_neg_1_14_port, Y(13) => 
                           out_shifter_neg_1_13_port, Y(12) => 
                           out_shifter_neg_1_12_port, Y(11) => 
                           out_shifter_neg_1_11_port, Y(10) => 
                           out_shifter_neg_1_10_port, Y(9) => 
                           out_shifter_neg_1_9_port, Y(8) => 
                           out_shifter_neg_1_8_port, Y(7) => 
                           out_shifter_neg_1_7_port, Y(6) => 
                           out_shifter_neg_1_6_port, Y(5) => 
                           out_shifter_neg_1_5_port, Y(4) => 
                           out_shifter_neg_1_4_port, Y(3) => 
                           out_shifter_neg_1_3_port, Y(2) => 
                           out_shifter_neg_1_2_port, Y(1) => 
                           out_shifter_neg_1_1_port, Y(0) => 
                           out_shifter_neg_1_0_port);
   COMP_2 : complementor_N16_6 port map( A(15) => out_shifter_2_15_port, A(14) 
                           => out_shifter_2_14_port, A(13) => 
                           out_shifter_2_13_port, A(12) => 
                           out_shifter_2_12_port, A(11) => 
                           out_shifter_2_11_port, A(10) => 
                           out_shifter_2_10_port, A(9) => out_shifter_2_9_port,
                           A(8) => out_shifter_2_8_port, A(7) => 
                           out_shifter_2_7_port, A(6) => out_shifter_2_6_port, 
                           A(5) => out_shifter_2_5_port, A(4) => 
                           out_shifter_2_4_port, A(3) => out_shifter_2_3_port, 
                           A(2) => out_shifter_2_2_port, A(1) => 
                           out_shifter_2_1_port, A(0) => out_shifter_2_0_port, 
                           Y(15) => out_shifter_neg_2_15_port, Y(14) => 
                           out_shifter_neg_2_14_port, Y(13) => 
                           out_shifter_neg_2_13_port, Y(12) => 
                           out_shifter_neg_2_12_port, Y(11) => 
                           out_shifter_neg_2_11_port, Y(10) => 
                           out_shifter_neg_2_10_port, Y(9) => 
                           out_shifter_neg_2_9_port, Y(8) => 
                           out_shifter_neg_2_8_port, Y(7) => 
                           out_shifter_neg_2_7_port, Y(6) => 
                           out_shifter_neg_2_6_port, Y(5) => 
                           out_shifter_neg_2_5_port, Y(4) => 
                           out_shifter_neg_2_4_port, Y(3) => 
                           out_shifter_neg_2_3_port, Y(2) => 
                           out_shifter_neg_2_2_port, Y(1) => 
                           out_shifter_neg_2_1_port, Y(0) => 
                           out_shifter_neg_2_0_port);
   COMP_3 : complementor_N16_5 port map( A(15) => out_shifter_3_15_port, A(14) 
                           => out_shifter_3_14_port, A(13) => 
                           out_shifter_3_13_port, A(12) => 
                           out_shifter_3_12_port, A(11) => 
                           out_shifter_3_11_port, A(10) => 
                           out_shifter_3_10_port, A(9) => out_shifter_3_9_port,
                           A(8) => out_shifter_3_8_port, A(7) => 
                           out_shifter_3_7_port, A(6) => out_shifter_3_6_port, 
                           A(5) => out_shifter_3_5_port, A(4) => 
                           out_shifter_3_4_port, A(3) => out_shifter_3_3_port, 
                           A(2) => out_shifter_3_2_port, A(1) => 
                           out_shifter_3_1_port, A(0) => out_shifter_3_0_port, 
                           Y(15) => out_shifter_neg_3_15_port, Y(14) => 
                           out_shifter_neg_3_14_port, Y(13) => 
                           out_shifter_neg_3_13_port, Y(12) => 
                           out_shifter_neg_3_12_port, Y(11) => 
                           out_shifter_neg_3_11_port, Y(10) => 
                           out_shifter_neg_3_10_port, Y(9) => 
                           out_shifter_neg_3_9_port, Y(8) => 
                           out_shifter_neg_3_8_port, Y(7) => 
                           out_shifter_neg_3_7_port, Y(6) => 
                           out_shifter_neg_3_6_port, Y(5) => 
                           out_shifter_neg_3_5_port, Y(4) => 
                           out_shifter_neg_3_4_port, Y(3) => 
                           out_shifter_neg_3_3_port, Y(2) => 
                           out_shifter_neg_3_2_port, Y(1) => 
                           out_shifter_neg_3_1_port, Y(0) => 
                           out_shifter_neg_3_0_port);
   COMP_4 : complementor_N16_4 port map( A(15) => out_shifter_4_15_port, A(14) 
                           => out_shifter_4_14_port, A(13) => 
                           out_shifter_4_13_port, A(12) => 
                           out_shifter_4_12_port, A(11) => 
                           out_shifter_4_11_port, A(10) => 
                           out_shifter_4_10_port, A(9) => out_shifter_4_9_port,
                           A(8) => out_shifter_4_8_port, A(7) => 
                           out_shifter_4_7_port, A(6) => out_shifter_4_6_port, 
                           A(5) => out_shifter_4_5_port, A(4) => 
                           out_shifter_4_4_port, A(3) => out_shifter_4_3_port, 
                           A(2) => out_shifter_4_2_port, A(1) => 
                           out_shifter_4_1_port, A(0) => out_shifter_4_0_port, 
                           Y(15) => out_shifter_neg_4_15_port, Y(14) => 
                           out_shifter_neg_4_14_port, Y(13) => 
                           out_shifter_neg_4_13_port, Y(12) => 
                           out_shifter_neg_4_12_port, Y(11) => 
                           out_shifter_neg_4_11_port, Y(10) => 
                           out_shifter_neg_4_10_port, Y(9) => 
                           out_shifter_neg_4_9_port, Y(8) => 
                           out_shifter_neg_4_8_port, Y(7) => 
                           out_shifter_neg_4_7_port, Y(6) => 
                           out_shifter_neg_4_6_port, Y(5) => 
                           out_shifter_neg_4_5_port, Y(4) => 
                           out_shifter_neg_4_4_port, Y(3) => 
                           out_shifter_neg_4_3_port, Y(2) => 
                           out_shifter_neg_4_2_port, Y(1) => 
                           out_shifter_neg_4_1_port, Y(0) => 
                           out_shifter_neg_4_0_port);
   COMP_5 : complementor_N16_3 port map( A(15) => out_shifter_5_15_port, A(14) 
                           => out_shifter_5_14_port, A(13) => 
                           out_shifter_5_13_port, A(12) => 
                           out_shifter_5_12_port, A(11) => 
                           out_shifter_5_11_port, A(10) => 
                           out_shifter_5_10_port, A(9) => out_shifter_5_9_port,
                           A(8) => out_shifter_5_8_port, A(7) => 
                           out_shifter_5_7_port, A(6) => out_shifter_5_6_port, 
                           A(5) => out_shifter_5_5_port, A(4) => 
                           out_shifter_5_4_port, A(3) => out_shifter_5_3_port, 
                           A(2) => out_shifter_5_2_port, A(1) => 
                           out_shifter_5_1_port, A(0) => out_shifter_5_0_port, 
                           Y(15) => out_shifter_neg_5_15_port, Y(14) => 
                           out_shifter_neg_5_14_port, Y(13) => 
                           out_shifter_neg_5_13_port, Y(12) => 
                           out_shifter_neg_5_12_port, Y(11) => 
                           out_shifter_neg_5_11_port, Y(10) => 
                           out_shifter_neg_5_10_port, Y(9) => 
                           out_shifter_neg_5_9_port, Y(8) => 
                           out_shifter_neg_5_8_port, Y(7) => 
                           out_shifter_neg_5_7_port, Y(6) => 
                           out_shifter_neg_5_6_port, Y(5) => 
                           out_shifter_neg_5_5_port, Y(4) => 
                           out_shifter_neg_5_4_port, Y(3) => 
                           out_shifter_neg_5_3_port, Y(2) => 
                           out_shifter_neg_5_2_port, Y(1) => 
                           out_shifter_neg_5_1_port, Y(0) => 
                           out_shifter_neg_5_0_port);
   COMP_6 : complementor_N16_2 port map( A(15) => out_shifter_6_15_port, A(14) 
                           => out_shifter_6_14_port, A(13) => 
                           out_shifter_6_13_port, A(12) => 
                           out_shifter_6_12_port, A(11) => 
                           out_shifter_6_11_port, A(10) => 
                           out_shifter_6_10_port, A(9) => out_shifter_6_9_port,
                           A(8) => out_shifter_6_8_port, A(7) => 
                           out_shifter_6_7_port, A(6) => out_shifter_6_6_port, 
                           A(5) => out_shifter_6_5_port, A(4) => 
                           out_shifter_6_4_port, A(3) => out_shifter_6_3_port, 
                           A(2) => out_shifter_6_2_port, A(1) => 
                           out_shifter_6_1_port, A(0) => out_shifter_6_0_port, 
                           Y(15) => out_shifter_neg_6_15_port, Y(14) => 
                           out_shifter_neg_6_14_port, Y(13) => 
                           out_shifter_neg_6_13_port, Y(12) => 
                           out_shifter_neg_6_12_port, Y(11) => 
                           out_shifter_neg_6_11_port, Y(10) => 
                           out_shifter_neg_6_10_port, Y(9) => 
                           out_shifter_neg_6_9_port, Y(8) => 
                           out_shifter_neg_6_8_port, Y(7) => 
                           out_shifter_neg_6_7_port, Y(6) => 
                           out_shifter_neg_6_6_port, Y(5) => 
                           out_shifter_neg_6_5_port, Y(4) => 
                           out_shifter_neg_6_4_port, Y(3) => 
                           out_shifter_neg_6_3_port, Y(2) => 
                           out_shifter_neg_6_2_port, Y(1) => 
                           out_shifter_neg_6_1_port, Y(0) => 
                           out_shifter_neg_6_0_port);
   COMP_7 : complementor_N16_1 port map( A(15) => out_shifter_7_15_port, A(14) 
                           => out_shifter_7_14_port, A(13) => 
                           out_shifter_7_13_port, A(12) => 
                           out_shifter_7_12_port, A(11) => 
                           out_shifter_7_11_port, A(10) => 
                           out_shifter_7_10_port, A(9) => out_shifter_7_9_port,
                           A(8) => out_shifter_7_8_port, A(7) => 
                           out_shifter_7_7_port, A(6) => out_shifter_7_6_port, 
                           A(5) => out_shifter_7_5_port, A(4) => 
                           out_shifter_7_4_port, A(3) => out_shifter_7_3_port, 
                           A(2) => out_shifter_7_2_port, A(1) => 
                           out_shifter_7_1_port, A(0) => out_shifter_7_0_port, 
                           Y(15) => out_shifter_neg_7_15_port, Y(14) => 
                           out_shifter_neg_7_14_port, Y(13) => 
                           out_shifter_neg_7_13_port, Y(12) => 
                           out_shifter_neg_7_12_port, Y(11) => 
                           out_shifter_neg_7_11_port, Y(10) => 
                           out_shifter_neg_7_10_port, Y(9) => 
                           out_shifter_neg_7_9_port, Y(8) => 
                           out_shifter_neg_7_8_port, Y(7) => 
                           out_shifter_neg_7_7_port, Y(6) => 
                           out_shifter_neg_7_6_port, Y(5) => 
                           out_shifter_neg_7_5_port, Y(4) => 
                           out_shifter_neg_7_4_port, Y(3) => 
                           out_shifter_neg_7_3_port, Y(2) => 
                           out_shifter_neg_7_2_port, Y(1) => 
                           out_shifter_neg_7_1_port, Y(0) => 
                           out_shifter_neg_7_0_port);
   MUX_0 : mux_8to1_N16_0 port map( A1(15) => X_Logic0_port, A1(14) => 
                           X_Logic0_port, A1(13) => X_Logic0_port, A1(12) => 
                           X_Logic0_port, A1(11) => X_Logic0_port, A1(10) => 
                           X_Logic0_port, A1(9) => X_Logic0_port, A1(8) => 
                           X_Logic0_port, A1(7) => X_Logic0_port, A1(6) => 
                           X_Logic0_port, A1(5) => X_Logic0_port, A1(4) => 
                           X_Logic0_port, A1(3) => X_Logic0_port, A1(2) => 
                           X_Logic0_port, A1(1) => X_Logic0_port, A1(0) => 
                           X_Logic0_port, A2(15) => out_shifter_0_15_port, 
                           A2(14) => out_shifter_0_14_port, A2(13) => 
                           out_shifter_0_13_port, A2(12) => 
                           out_shifter_0_12_port, A2(11) => 
                           out_shifter_0_11_port, A2(10) => 
                           out_shifter_0_10_port, A2(9) => out_shifter_0_9_port
                           , A2(8) => out_shifter_0_8_port, A2(7) => 
                           out_shifter_0_7_port, A2(6) => out_shifter_0_6_port,
                           A2(5) => out_shifter_0_5_port, A2(4) => 
                           out_shifter_0_4_port, A2(3) => out_shifter_0_3_port,
                           A2(2) => out_shifter_0_2_port, A2(1) => 
                           out_shifter_0_1_port, A2(0) => out_shifter_0_0_port,
                           A3(15) => out_shifter_0_15_port, A3(14) => 
                           out_shifter_0_14_port, A3(13) => 
                           out_shifter_0_13_port, A3(12) => 
                           out_shifter_0_12_port, A3(11) => 
                           out_shifter_0_11_port, A3(10) => 
                           out_shifter_0_10_port, A3(9) => out_shifter_0_9_port
                           , A3(8) => out_shifter_0_8_port, A3(7) => 
                           out_shifter_0_7_port, A3(6) => out_shifter_0_6_port,
                           A3(5) => out_shifter_0_5_port, A3(4) => 
                           out_shifter_0_4_port, A3(3) => out_shifter_0_3_port,
                           A3(2) => out_shifter_0_2_port, A3(1) => 
                           out_shifter_0_1_port, A3(0) => out_shifter_0_0_port,
                           A4(15) => out_shifter_1_15_port, A4(14) => 
                           out_shifter_1_14_port, A4(13) => 
                           out_shifter_1_13_port, A4(12) => 
                           out_shifter_1_12_port, A4(11) => 
                           out_shifter_1_11_port, A4(10) => 
                           out_shifter_1_10_port, A4(9) => out_shifter_1_9_port
                           , A4(8) => out_shifter_1_8_port, A4(7) => 
                           out_shifter_1_7_port, A4(6) => out_shifter_1_6_port,
                           A4(5) => out_shifter_1_5_port, A4(4) => 
                           out_shifter_1_4_port, A4(3) => out_shifter_1_3_port,
                           A4(2) => out_shifter_1_2_port, A4(1) => 
                           out_shifter_1_1_port, A4(0) => out_shifter_1_0_port,
                           A5(15) => out_shifter_neg_1_15_port, A5(14) => 
                           out_shifter_neg_1_14_port, A5(13) => 
                           out_shifter_neg_1_13_port, A5(12) => 
                           out_shifter_neg_1_12_port, A5(11) => 
                           out_shifter_neg_1_11_port, A5(10) => 
                           out_shifter_neg_1_10_port, A5(9) => 
                           out_shifter_neg_1_9_port, A5(8) => 
                           out_shifter_neg_1_8_port, A5(7) => 
                           out_shifter_neg_1_7_port, A5(6) => 
                           out_shifter_neg_1_6_port, A5(5) => 
                           out_shifter_neg_1_5_port, A5(4) => 
                           out_shifter_neg_1_4_port, A5(3) => 
                           out_shifter_neg_1_3_port, A5(2) => 
                           out_shifter_neg_1_2_port, A5(1) => 
                           out_shifter_neg_1_1_port, A5(0) => 
                           out_shifter_neg_1_0_port, A6(15) => 
                           out_shifter_neg_0_15_port, A6(14) => 
                           out_shifter_neg_0_14_port, A6(13) => 
                           out_shifter_neg_0_13_port, A6(12) => 
                           out_shifter_neg_0_12_port, A6(11) => 
                           out_shifter_neg_0_11_port, A6(10) => 
                           out_shifter_neg_0_10_port, A6(9) => 
                           out_shifter_neg_0_9_port, A6(8) => 
                           out_shifter_neg_0_8_port, A6(7) => 
                           out_shifter_neg_0_7_port, A6(6) => 
                           out_shifter_neg_0_6_port, A6(5) => 
                           out_shifter_neg_0_5_port, A6(4) => 
                           out_shifter_neg_0_4_port, A6(3) => 
                           out_shifter_neg_0_3_port, A6(2) => 
                           out_shifter_neg_0_2_port, A6(1) => 
                           out_shifter_neg_0_1_port, A6(0) => 
                           out_shifter_neg_0_0_port, A7(15) => 
                           out_shifter_neg_0_15_port, A7(14) => 
                           out_shifter_neg_0_14_port, A7(13) => 
                           out_shifter_neg_0_13_port, A7(12) => 
                           out_shifter_neg_0_12_port, A7(11) => 
                           out_shifter_neg_0_11_port, A7(10) => 
                           out_shifter_neg_0_10_port, A7(9) => 
                           out_shifter_neg_0_9_port, A7(8) => 
                           out_shifter_neg_0_8_port, A7(7) => 
                           out_shifter_neg_0_7_port, A7(6) => 
                           out_shifter_neg_0_6_port, A7(5) => 
                           out_shifter_neg_0_5_port, A7(4) => 
                           out_shifter_neg_0_4_port, A7(3) => 
                           out_shifter_neg_0_3_port, A7(2) => 
                           out_shifter_neg_0_2_port, A7(1) => 
                           out_shifter_neg_0_1_port, A7(0) => 
                           out_shifter_neg_0_0_port, A8(15) => X_Logic0_port, 
                           A8(14) => X_Logic0_port, A8(13) => X_Logic0_port, 
                           A8(12) => X_Logic0_port, A8(11) => X_Logic0_port, 
                           A8(10) => X_Logic0_port, A8(9) => X_Logic0_port, 
                           A8(8) => X_Logic0_port, A8(7) => X_Logic0_port, 
                           A8(6) => X_Logic0_port, A8(5) => X_Logic0_port, 
                           A8(4) => X_Logic0_port, A8(3) => X_Logic0_port, 
                           A8(2) => X_Logic0_port, A8(1) => X_Logic0_port, 
                           A8(0) => X_Logic0_port, S(2) => sel_muxes_2_port, 
                           S(1) => sel_muxes_1_port, S(0) => sel_muxes_0_port, 
                           Y(15) => out_muxes_0_15_port, Y(14) => 
                           out_muxes_0_14_port, Y(13) => out_muxes_0_13_port, 
                           Y(12) => out_muxes_0_12_port, Y(11) => 
                           out_muxes_0_11_port, Y(10) => out_muxes_0_10_port, 
                           Y(9) => out_muxes_0_9_port, Y(8) => 
                           out_muxes_0_8_port, Y(7) => out_muxes_0_7_port, Y(6)
                           => out_muxes_0_6_port, Y(5) => out_muxes_0_5_port, 
                           Y(4) => out_muxes_0_4_port, Y(3) => 
                           out_muxes_0_3_port, Y(2) => out_muxes_0_2_port, Y(1)
                           => out_muxes_0_1_port, Y(0) => out_muxes_0_0_port);
   MUX_1 : mux_8to1_N16_3 port map( A1(15) => X_Logic0_port, A1(14) => 
                           X_Logic0_port, A1(13) => X_Logic0_port, A1(12) => 
                           X_Logic0_port, A1(11) => X_Logic0_port, A1(10) => 
                           X_Logic0_port, A1(9) => X_Logic0_port, A1(8) => 
                           X_Logic0_port, A1(7) => X_Logic0_port, A1(6) => 
                           X_Logic0_port, A1(5) => X_Logic0_port, A1(4) => 
                           X_Logic0_port, A1(3) => X_Logic0_port, A1(2) => 
                           X_Logic0_port, A1(1) => X_Logic0_port, A1(0) => 
                           X_Logic0_port, A2(15) => out_shifter_2_15_port, 
                           A2(14) => out_shifter_2_14_port, A2(13) => 
                           out_shifter_2_13_port, A2(12) => 
                           out_shifter_2_12_port, A2(11) => 
                           out_shifter_2_11_port, A2(10) => 
                           out_shifter_2_10_port, A2(9) => out_shifter_2_9_port
                           , A2(8) => out_shifter_2_8_port, A2(7) => 
                           out_shifter_2_7_port, A2(6) => out_shifter_2_6_port,
                           A2(5) => out_shifter_2_5_port, A2(4) => 
                           out_shifter_2_4_port, A2(3) => out_shifter_2_3_port,
                           A2(2) => out_shifter_2_2_port, A2(1) => 
                           out_shifter_2_1_port, A2(0) => out_shifter_2_0_port,
                           A3(15) => out_shifter_2_15_port, A3(14) => 
                           out_shifter_2_14_port, A3(13) => 
                           out_shifter_2_13_port, A3(12) => 
                           out_shifter_2_12_port, A3(11) => 
                           out_shifter_2_11_port, A3(10) => 
                           out_shifter_2_10_port, A3(9) => out_shifter_2_9_port
                           , A3(8) => out_shifter_2_8_port, A3(7) => 
                           out_shifter_2_7_port, A3(6) => out_shifter_2_6_port,
                           A3(5) => out_shifter_2_5_port, A3(4) => 
                           out_shifter_2_4_port, A3(3) => out_shifter_2_3_port,
                           A3(2) => out_shifter_2_2_port, A3(1) => 
                           out_shifter_2_1_port, A3(0) => out_shifter_2_0_port,
                           A4(15) => out_shifter_3_15_port, A4(14) => 
                           out_shifter_3_14_port, A4(13) => 
                           out_shifter_3_13_port, A4(12) => 
                           out_shifter_3_12_port, A4(11) => 
                           out_shifter_3_11_port, A4(10) => 
                           out_shifter_3_10_port, A4(9) => out_shifter_3_9_port
                           , A4(8) => out_shifter_3_8_port, A4(7) => 
                           out_shifter_3_7_port, A4(6) => out_shifter_3_6_port,
                           A4(5) => out_shifter_3_5_port, A4(4) => 
                           out_shifter_3_4_port, A4(3) => out_shifter_3_3_port,
                           A4(2) => out_shifter_3_2_port, A4(1) => 
                           out_shifter_3_1_port, A4(0) => out_shifter_3_0_port,
                           A5(15) => out_shifter_neg_3_15_port, A5(14) => 
                           out_shifter_neg_3_14_port, A5(13) => 
                           out_shifter_neg_3_13_port, A5(12) => 
                           out_shifter_neg_3_12_port, A5(11) => 
                           out_shifter_neg_3_11_port, A5(10) => 
                           out_shifter_neg_3_10_port, A5(9) => 
                           out_shifter_neg_3_9_port, A5(8) => 
                           out_shifter_neg_3_8_port, A5(7) => 
                           out_shifter_neg_3_7_port, A5(6) => 
                           out_shifter_neg_3_6_port, A5(5) => 
                           out_shifter_neg_3_5_port, A5(4) => 
                           out_shifter_neg_3_4_port, A5(3) => 
                           out_shifter_neg_3_3_port, A5(2) => 
                           out_shifter_neg_3_2_port, A5(1) => 
                           out_shifter_neg_3_1_port, A5(0) => 
                           out_shifter_neg_3_0_port, A6(15) => 
                           out_shifter_neg_2_15_port, A6(14) => 
                           out_shifter_neg_2_14_port, A6(13) => 
                           out_shifter_neg_2_13_port, A6(12) => 
                           out_shifter_neg_2_12_port, A6(11) => 
                           out_shifter_neg_2_11_port, A6(10) => 
                           out_shifter_neg_2_10_port, A6(9) => 
                           out_shifter_neg_2_9_port, A6(8) => 
                           out_shifter_neg_2_8_port, A6(7) => 
                           out_shifter_neg_2_7_port, A6(6) => 
                           out_shifter_neg_2_6_port, A6(5) => 
                           out_shifter_neg_2_5_port, A6(4) => 
                           out_shifter_neg_2_4_port, A6(3) => 
                           out_shifter_neg_2_3_port, A6(2) => 
                           out_shifter_neg_2_2_port, A6(1) => 
                           out_shifter_neg_2_1_port, A6(0) => 
                           out_shifter_neg_2_0_port, A7(15) => 
                           out_shifter_neg_2_15_port, A7(14) => 
                           out_shifter_neg_2_14_port, A7(13) => 
                           out_shifter_neg_2_13_port, A7(12) => 
                           out_shifter_neg_2_12_port, A7(11) => 
                           out_shifter_neg_2_11_port, A7(10) => 
                           out_shifter_neg_2_10_port, A7(9) => 
                           out_shifter_neg_2_9_port, A7(8) => 
                           out_shifter_neg_2_8_port, A7(7) => 
                           out_shifter_neg_2_7_port, A7(6) => 
                           out_shifter_neg_2_6_port, A7(5) => 
                           out_shifter_neg_2_5_port, A7(4) => 
                           out_shifter_neg_2_4_port, A7(3) => 
                           out_shifter_neg_2_3_port, A7(2) => 
                           out_shifter_neg_2_2_port, A7(1) => 
                           out_shifter_neg_2_1_port, A7(0) => 
                           out_shifter_neg_2_0_port, A8(15) => X_Logic0_port, 
                           A8(14) => X_Logic0_port, A8(13) => X_Logic0_port, 
                           A8(12) => X_Logic0_port, A8(11) => X_Logic0_port, 
                           A8(10) => X_Logic0_port, A8(9) => X_Logic0_port, 
                           A8(8) => X_Logic0_port, A8(7) => X_Logic0_port, 
                           A8(6) => X_Logic0_port, A8(5) => X_Logic0_port, 
                           A8(4) => X_Logic0_port, A8(3) => X_Logic0_port, 
                           A8(2) => X_Logic0_port, A8(1) => X_Logic0_port, 
                           A8(0) => X_Logic0_port, S(2) => sel_muxes_5_port, 
                           S(1) => sel_muxes_4_port, S(0) => sel_muxes_3_port, 
                           Y(15) => out_muxes_1_15_port, Y(14) => 
                           out_muxes_1_14_port, Y(13) => out_muxes_1_13_port, 
                           Y(12) => out_muxes_1_12_port, Y(11) => 
                           out_muxes_1_11_port, Y(10) => out_muxes_1_10_port, 
                           Y(9) => out_muxes_1_9_port, Y(8) => 
                           out_muxes_1_8_port, Y(7) => out_muxes_1_7_port, Y(6)
                           => out_muxes_1_6_port, Y(5) => out_muxes_1_5_port, 
                           Y(4) => out_muxes_1_4_port, Y(3) => 
                           out_muxes_1_3_port, Y(2) => out_muxes_1_2_port, Y(1)
                           => out_muxes_1_1_port, Y(0) => out_muxes_1_0_port);
   MUX_2 : mux_8to1_N16_2 port map( A1(15) => X_Logic0_port, A1(14) => 
                           X_Logic0_port, A1(13) => X_Logic0_port, A1(12) => 
                           X_Logic0_port, A1(11) => X_Logic0_port, A1(10) => 
                           X_Logic0_port, A1(9) => X_Logic0_port, A1(8) => 
                           X_Logic0_port, A1(7) => X_Logic0_port, A1(6) => 
                           X_Logic0_port, A1(5) => X_Logic0_port, A1(4) => 
                           X_Logic0_port, A1(3) => X_Logic0_port, A1(2) => 
                           X_Logic0_port, A1(1) => X_Logic0_port, A1(0) => 
                           X_Logic0_port, A2(15) => out_shifter_4_15_port, 
                           A2(14) => out_shifter_4_14_port, A2(13) => 
                           out_shifter_4_13_port, A2(12) => 
                           out_shifter_4_12_port, A2(11) => 
                           out_shifter_4_11_port, A2(10) => 
                           out_shifter_4_10_port, A2(9) => out_shifter_4_9_port
                           , A2(8) => out_shifter_4_8_port, A2(7) => 
                           out_shifter_4_7_port, A2(6) => out_shifter_4_6_port,
                           A2(5) => out_shifter_4_5_port, A2(4) => 
                           out_shifter_4_4_port, A2(3) => out_shifter_4_3_port,
                           A2(2) => out_shifter_4_2_port, A2(1) => 
                           out_shifter_4_1_port, A2(0) => out_shifter_4_0_port,
                           A3(15) => out_shifter_4_15_port, A3(14) => 
                           out_shifter_4_14_port, A3(13) => 
                           out_shifter_4_13_port, A3(12) => 
                           out_shifter_4_12_port, A3(11) => 
                           out_shifter_4_11_port, A3(10) => 
                           out_shifter_4_10_port, A3(9) => out_shifter_4_9_port
                           , A3(8) => out_shifter_4_8_port, A3(7) => 
                           out_shifter_4_7_port, A3(6) => out_shifter_4_6_port,
                           A3(5) => out_shifter_4_5_port, A3(4) => 
                           out_shifter_4_4_port, A3(3) => out_shifter_4_3_port,
                           A3(2) => out_shifter_4_2_port, A3(1) => 
                           out_shifter_4_1_port, A3(0) => out_shifter_4_0_port,
                           A4(15) => out_shifter_5_15_port, A4(14) => 
                           out_shifter_5_14_port, A4(13) => 
                           out_shifter_5_13_port, A4(12) => 
                           out_shifter_5_12_port, A4(11) => 
                           out_shifter_5_11_port, A4(10) => 
                           out_shifter_5_10_port, A4(9) => out_shifter_5_9_port
                           , A4(8) => out_shifter_5_8_port, A4(7) => 
                           out_shifter_5_7_port, A4(6) => out_shifter_5_6_port,
                           A4(5) => out_shifter_5_5_port, A4(4) => 
                           out_shifter_5_4_port, A4(3) => out_shifter_5_3_port,
                           A4(2) => out_shifter_5_2_port, A4(1) => 
                           out_shifter_5_1_port, A4(0) => out_shifter_5_0_port,
                           A5(15) => out_shifter_neg_5_15_port, A5(14) => 
                           out_shifter_neg_5_14_port, A5(13) => 
                           out_shifter_neg_5_13_port, A5(12) => 
                           out_shifter_neg_5_12_port, A5(11) => 
                           out_shifter_neg_5_11_port, A5(10) => 
                           out_shifter_neg_5_10_port, A5(9) => 
                           out_shifter_neg_5_9_port, A5(8) => 
                           out_shifter_neg_5_8_port, A5(7) => 
                           out_shifter_neg_5_7_port, A5(6) => 
                           out_shifter_neg_5_6_port, A5(5) => 
                           out_shifter_neg_5_5_port, A5(4) => 
                           out_shifter_neg_5_4_port, A5(3) => 
                           out_shifter_neg_5_3_port, A5(2) => 
                           out_shifter_neg_5_2_port, A5(1) => 
                           out_shifter_neg_5_1_port, A5(0) => 
                           out_shifter_neg_5_0_port, A6(15) => 
                           out_shifter_neg_4_15_port, A6(14) => 
                           out_shifter_neg_4_14_port, A6(13) => 
                           out_shifter_neg_4_13_port, A6(12) => 
                           out_shifter_neg_4_12_port, A6(11) => 
                           out_shifter_neg_4_11_port, A6(10) => 
                           out_shifter_neg_4_10_port, A6(9) => 
                           out_shifter_neg_4_9_port, A6(8) => 
                           out_shifter_neg_4_8_port, A6(7) => 
                           out_shifter_neg_4_7_port, A6(6) => 
                           out_shifter_neg_4_6_port, A6(5) => 
                           out_shifter_neg_4_5_port, A6(4) => 
                           out_shifter_neg_4_4_port, A6(3) => 
                           out_shifter_neg_4_3_port, A6(2) => 
                           out_shifter_neg_4_2_port, A6(1) => 
                           out_shifter_neg_4_1_port, A6(0) => 
                           out_shifter_neg_4_0_port, A7(15) => 
                           out_shifter_neg_4_15_port, A7(14) => 
                           out_shifter_neg_4_14_port, A7(13) => 
                           out_shifter_neg_4_13_port, A7(12) => 
                           out_shifter_neg_4_12_port, A7(11) => 
                           out_shifter_neg_4_11_port, A7(10) => 
                           out_shifter_neg_4_10_port, A7(9) => 
                           out_shifter_neg_4_9_port, A7(8) => 
                           out_shifter_neg_4_8_port, A7(7) => 
                           out_shifter_neg_4_7_port, A7(6) => 
                           out_shifter_neg_4_6_port, A7(5) => 
                           out_shifter_neg_4_5_port, A7(4) => 
                           out_shifter_neg_4_4_port, A7(3) => 
                           out_shifter_neg_4_3_port, A7(2) => 
                           out_shifter_neg_4_2_port, A7(1) => 
                           out_shifter_neg_4_1_port, A7(0) => 
                           out_shifter_neg_4_0_port, A8(15) => X_Logic0_port, 
                           A8(14) => X_Logic0_port, A8(13) => X_Logic0_port, 
                           A8(12) => X_Logic0_port, A8(11) => X_Logic0_port, 
                           A8(10) => X_Logic0_port, A8(9) => X_Logic0_port, 
                           A8(8) => X_Logic0_port, A8(7) => X_Logic0_port, 
                           A8(6) => X_Logic0_port, A8(5) => X_Logic0_port, 
                           A8(4) => X_Logic0_port, A8(3) => X_Logic0_port, 
                           A8(2) => X_Logic0_port, A8(1) => X_Logic0_port, 
                           A8(0) => X_Logic0_port, S(2) => sel_muxes_8_port, 
                           S(1) => sel_muxes_7_port, S(0) => sel_muxes_6_port, 
                           Y(15) => out_muxes_2_15_port, Y(14) => 
                           out_muxes_2_14_port, Y(13) => out_muxes_2_13_port, 
                           Y(12) => out_muxes_2_12_port, Y(11) => 
                           out_muxes_2_11_port, Y(10) => out_muxes_2_10_port, 
                           Y(9) => out_muxes_2_9_port, Y(8) => 
                           out_muxes_2_8_port, Y(7) => out_muxes_2_7_port, Y(6)
                           => out_muxes_2_6_port, Y(5) => out_muxes_2_5_port, 
                           Y(4) => out_muxes_2_4_port, Y(3) => 
                           out_muxes_2_3_port, Y(2) => out_muxes_2_2_port, Y(1)
                           => out_muxes_2_1_port, Y(0) => out_muxes_2_0_port);
   MUX_3 : mux_8to1_N16_1 port map( A1(15) => X_Logic0_port, A1(14) => 
                           X_Logic0_port, A1(13) => X_Logic0_port, A1(12) => 
                           X_Logic0_port, A1(11) => X_Logic0_port, A1(10) => 
                           X_Logic0_port, A1(9) => X_Logic0_port, A1(8) => 
                           X_Logic0_port, A1(7) => X_Logic0_port, A1(6) => 
                           X_Logic0_port, A1(5) => X_Logic0_port, A1(4) => 
                           X_Logic0_port, A1(3) => X_Logic0_port, A1(2) => 
                           X_Logic0_port, A1(1) => X_Logic0_port, A1(0) => 
                           X_Logic0_port, A2(15) => out_shifter_6_15_port, 
                           A2(14) => out_shifter_6_14_port, A2(13) => 
                           out_shifter_6_13_port, A2(12) => 
                           out_shifter_6_12_port, A2(11) => 
                           out_shifter_6_11_port, A2(10) => 
                           out_shifter_6_10_port, A2(9) => out_shifter_6_9_port
                           , A2(8) => out_shifter_6_8_port, A2(7) => 
                           out_shifter_6_7_port, A2(6) => out_shifter_6_6_port,
                           A2(5) => out_shifter_6_5_port, A2(4) => 
                           out_shifter_6_4_port, A2(3) => out_shifter_6_3_port,
                           A2(2) => out_shifter_6_2_port, A2(1) => 
                           out_shifter_6_1_port, A2(0) => out_shifter_6_0_port,
                           A3(15) => out_shifter_6_15_port, A3(14) => 
                           out_shifter_6_14_port, A3(13) => 
                           out_shifter_6_13_port, A3(12) => 
                           out_shifter_6_12_port, A3(11) => 
                           out_shifter_6_11_port, A3(10) => 
                           out_shifter_6_10_port, A3(9) => out_shifter_6_9_port
                           , A3(8) => out_shifter_6_8_port, A3(7) => 
                           out_shifter_6_7_port, A3(6) => out_shifter_6_6_port,
                           A3(5) => out_shifter_6_5_port, A3(4) => 
                           out_shifter_6_4_port, A3(3) => out_shifter_6_3_port,
                           A3(2) => out_shifter_6_2_port, A3(1) => 
                           out_shifter_6_1_port, A3(0) => out_shifter_6_0_port,
                           A4(15) => out_shifter_7_15_port, A4(14) => 
                           out_shifter_7_14_port, A4(13) => 
                           out_shifter_7_13_port, A4(12) => 
                           out_shifter_7_12_port, A4(11) => 
                           out_shifter_7_11_port, A4(10) => 
                           out_shifter_7_10_port, A4(9) => out_shifter_7_9_port
                           , A4(8) => out_shifter_7_8_port, A4(7) => 
                           out_shifter_7_7_port, A4(6) => out_shifter_7_6_port,
                           A4(5) => out_shifter_7_5_port, A4(4) => 
                           out_shifter_7_4_port, A4(3) => out_shifter_7_3_port,
                           A4(2) => out_shifter_7_2_port, A4(1) => 
                           out_shifter_7_1_port, A4(0) => out_shifter_7_0_port,
                           A5(15) => out_shifter_neg_7_15_port, A5(14) => 
                           out_shifter_neg_7_14_port, A5(13) => 
                           out_shifter_neg_7_13_port, A5(12) => 
                           out_shifter_neg_7_12_port, A5(11) => 
                           out_shifter_neg_7_11_port, A5(10) => 
                           out_shifter_neg_7_10_port, A5(9) => 
                           out_shifter_neg_7_9_port, A5(8) => 
                           out_shifter_neg_7_8_port, A5(7) => 
                           out_shifter_neg_7_7_port, A5(6) => 
                           out_shifter_neg_7_6_port, A5(5) => 
                           out_shifter_neg_7_5_port, A5(4) => 
                           out_shifter_neg_7_4_port, A5(3) => 
                           out_shifter_neg_7_3_port, A5(2) => 
                           out_shifter_neg_7_2_port, A5(1) => 
                           out_shifter_neg_7_1_port, A5(0) => 
                           out_shifter_neg_7_0_port, A6(15) => 
                           out_shifter_neg_6_15_port, A6(14) => 
                           out_shifter_neg_6_14_port, A6(13) => 
                           out_shifter_neg_6_13_port, A6(12) => 
                           out_shifter_neg_6_12_port, A6(11) => 
                           out_shifter_neg_6_11_port, A6(10) => 
                           out_shifter_neg_6_10_port, A6(9) => 
                           out_shifter_neg_6_9_port, A6(8) => 
                           out_shifter_neg_6_8_port, A6(7) => 
                           out_shifter_neg_6_7_port, A6(6) => 
                           out_shifter_neg_6_6_port, A6(5) => 
                           out_shifter_neg_6_5_port, A6(4) => 
                           out_shifter_neg_6_4_port, A6(3) => 
                           out_shifter_neg_6_3_port, A6(2) => 
                           out_shifter_neg_6_2_port, A6(1) => 
                           out_shifter_neg_6_1_port, A6(0) => 
                           out_shifter_neg_6_0_port, A7(15) => 
                           out_shifter_neg_6_15_port, A7(14) => 
                           out_shifter_neg_6_14_port, A7(13) => 
                           out_shifter_neg_6_13_port, A7(12) => 
                           out_shifter_neg_6_12_port, A7(11) => 
                           out_shifter_neg_6_11_port, A7(10) => 
                           out_shifter_neg_6_10_port, A7(9) => 
                           out_shifter_neg_6_9_port, A7(8) => 
                           out_shifter_neg_6_8_port, A7(7) => 
                           out_shifter_neg_6_7_port, A7(6) => 
                           out_shifter_neg_6_6_port, A7(5) => 
                           out_shifter_neg_6_5_port, A7(4) => 
                           out_shifter_neg_6_4_port, A7(3) => 
                           out_shifter_neg_6_3_port, A7(2) => 
                           out_shifter_neg_6_2_port, A7(1) => 
                           out_shifter_neg_6_1_port, A7(0) => 
                           out_shifter_neg_6_0_port, A8(15) => X_Logic0_port, 
                           A8(14) => X_Logic0_port, A8(13) => X_Logic0_port, 
                           A8(12) => X_Logic0_port, A8(11) => X_Logic0_port, 
                           A8(10) => X_Logic0_port, A8(9) => X_Logic0_port, 
                           A8(8) => X_Logic0_port, A8(7) => X_Logic0_port, 
                           A8(6) => X_Logic0_port, A8(5) => X_Logic0_port, 
                           A8(4) => X_Logic0_port, A8(3) => X_Logic0_port, 
                           A8(2) => X_Logic0_port, A8(1) => X_Logic0_port, 
                           A8(0) => X_Logic0_port, S(2) => sel_muxes_11_port, 
                           S(1) => sel_muxes_10_port, S(0) => sel_muxes_9_port,
                           Y(15) => out_muxes_3_15_port, Y(14) => 
                           out_muxes_3_14_port, Y(13) => out_muxes_3_13_port, 
                           Y(12) => out_muxes_3_12_port, Y(11) => 
                           out_muxes_3_11_port, Y(10) => out_muxes_3_10_port, 
                           Y(9) => out_muxes_3_9_port, Y(8) => 
                           out_muxes_3_8_port, Y(7) => out_muxes_3_7_port, Y(6)
                           => out_muxes_3_6_port, Y(5) => out_muxes_3_5_port, 
                           Y(4) => out_muxes_3_4_port, Y(3) => 
                           out_muxes_3_3_port, Y(2) => out_muxes_3_2_port, Y(1)
                           => out_muxes_3_1_port, Y(0) => out_muxes_3_0_port);
   SUM0_0 : P4_adder_N16_Nbit_blocks4_0 port map( A(15) => out_muxes_0_15_port,
                           A(14) => out_muxes_0_14_port, A(13) => 
                           out_muxes_0_13_port, A(12) => out_muxes_0_12_port, 
                           A(11) => out_muxes_0_11_port, A(10) => 
                           out_muxes_0_10_port, A(9) => out_muxes_0_9_port, 
                           A(8) => out_muxes_0_8_port, A(7) => 
                           out_muxes_0_7_port, A(6) => out_muxes_0_6_port, A(5)
                           => out_muxes_0_5_port, A(4) => out_muxes_0_4_port, 
                           A(3) => out_muxes_0_3_port, A(2) => 
                           out_muxes_0_2_port, A(1) => out_muxes_0_1_port, A(0)
                           => out_muxes_0_0_port, B(15) => out_muxes_1_15_port,
                           B(14) => out_muxes_1_14_port, B(13) => 
                           out_muxes_1_13_port, B(12) => out_muxes_1_12_port, 
                           B(11) => out_muxes_1_11_port, B(10) => 
                           out_muxes_1_10_port, B(9) => out_muxes_1_9_port, 
                           B(8) => out_muxes_1_8_port, B(7) => 
                           out_muxes_1_7_port, B(6) => out_muxes_1_6_port, B(5)
                           => out_muxes_1_5_port, B(4) => out_muxes_1_4_port, 
                           B(3) => out_muxes_1_3_port, B(2) => 
                           out_muxes_1_2_port, B(1) => out_muxes_1_1_port, B(0)
                           => out_muxes_1_0_port, Cin => X_Logic0_port, S(15) 
                           => out_adder_0_15_port, S(14) => out_adder_0_14_port
                           , S(13) => out_adder_0_13_port, S(12) => 
                           out_adder_0_12_port, S(11) => out_adder_0_11_port, 
                           S(10) => out_adder_0_10_port, S(9) => 
                           out_adder_0_9_port, S(8) => out_adder_0_8_port, S(7)
                           => out_adder_0_7_port, S(6) => out_adder_0_6_port, 
                           S(5) => out_adder_0_5_port, S(4) => 
                           out_adder_0_4_port, S(3) => out_adder_0_3_port, S(2)
                           => out_adder_0_2_port, S(1) => out_adder_0_1_port, 
                           S(0) => out_adder_0_0_port, Cout => n_1123);
   SUMn_1 : P4_adder_N16_Nbit_blocks4_2 port map( A(15) => out_muxes_2_15_port,
                           A(14) => out_muxes_2_14_port, A(13) => 
                           out_muxes_2_13_port, A(12) => out_muxes_2_12_port, 
                           A(11) => out_muxes_2_11_port, A(10) => 
                           out_muxes_2_10_port, A(9) => out_muxes_2_9_port, 
                           A(8) => out_muxes_2_8_port, A(7) => 
                           out_muxes_2_7_port, A(6) => out_muxes_2_6_port, A(5)
                           => out_muxes_2_5_port, A(4) => out_muxes_2_4_port, 
                           A(3) => out_muxes_2_3_port, A(2) => 
                           out_muxes_2_2_port, A(1) => out_muxes_2_1_port, A(0)
                           => out_muxes_2_0_port, B(15) => out_adder_0_15_port,
                           B(14) => out_adder_0_14_port, B(13) => 
                           out_adder_0_13_port, B(12) => out_adder_0_12_port, 
                           B(11) => out_adder_0_11_port, B(10) => 
                           out_adder_0_10_port, B(9) => out_adder_0_9_port, 
                           B(8) => out_adder_0_8_port, B(7) => 
                           out_adder_0_7_port, B(6) => out_adder_0_6_port, B(5)
                           => out_adder_0_5_port, B(4) => out_adder_0_4_port, 
                           B(3) => out_adder_0_3_port, B(2) => 
                           out_adder_0_2_port, B(1) => out_adder_0_1_port, B(0)
                           => out_adder_0_0_port, Cin => X_Logic0_port, S(15) 
                           => out_adder_1_15_port, S(14) => out_adder_1_14_port
                           , S(13) => out_adder_1_13_port, S(12) => 
                           out_adder_1_12_port, S(11) => out_adder_1_11_port, 
                           S(10) => out_adder_1_10_port, S(9) => 
                           out_adder_1_9_port, S(8) => out_adder_1_8_port, S(7)
                           => out_adder_1_7_port, S(6) => out_adder_1_6_port, 
                           S(5) => out_adder_1_5_port, S(4) => 
                           out_adder_1_4_port, S(3) => out_adder_1_3_port, S(2)
                           => out_adder_1_2_port, S(1) => out_adder_1_1_port, 
                           S(0) => out_adder_1_0_port, Cout => n_1124);
   SUMn_2 : P4_adder_N16_Nbit_blocks4_1 port map( A(15) => out_muxes_3_15_port,
                           A(14) => out_muxes_3_14_port, A(13) => 
                           out_muxes_3_13_port, A(12) => out_muxes_3_12_port, 
                           A(11) => out_muxes_3_11_port, A(10) => 
                           out_muxes_3_10_port, A(9) => out_muxes_3_9_port, 
                           A(8) => out_muxes_3_8_port, A(7) => 
                           out_muxes_3_7_port, A(6) => out_muxes_3_6_port, A(5)
                           => out_muxes_3_5_port, A(4) => out_muxes_3_4_port, 
                           A(3) => out_muxes_3_3_port, A(2) => 
                           out_muxes_3_2_port, A(1) => out_muxes_3_1_port, A(0)
                           => out_muxes_3_0_port, B(15) => out_adder_1_15_port,
                           B(14) => out_adder_1_14_port, B(13) => 
                           out_adder_1_13_port, B(12) => out_adder_1_12_port, 
                           B(11) => out_adder_1_11_port, B(10) => 
                           out_adder_1_10_port, B(9) => out_adder_1_9_port, 
                           B(8) => out_adder_1_8_port, B(7) => 
                           out_adder_1_7_port, B(6) => out_adder_1_6_port, B(5)
                           => out_adder_1_5_port, B(4) => out_adder_1_4_port, 
                           B(3) => out_adder_1_3_port, B(2) => 
                           out_adder_1_2_port, B(1) => out_adder_1_1_port, B(0)
                           => out_adder_1_0_port, Cin => X_Logic0_port, S(15) 
                           => Y(15), S(14) => Y(14), S(13) => Y(13), S(12) => 
                           Y(12), S(11) => Y(11), S(10) => Y(10), S(9) => Y(9),
                           S(8) => Y(8), S(7) => Y(7), S(6) => Y(6), S(5) => 
                           Y(5), S(4) => Y(4), S(3) => Y(3), S(2) => Y(2), S(1)
                           => Y(1), S(0) => Y(0), Cout => n_1125);

end SYN_ARCHSTRUCT;
